// DE2_115_QSYS.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module DE2_115_QSYS (
		input  wire [7:0]  camera_blue_in_external_connection_export,  //  camera_blue_in_external_connection.export
		input  wire [7:0]  camera_green_in_external_connection_export, // camera_green_in_external_connection.export
		input  wire [7:0]  camera_red_in_external_connection_export,   //   camera_red_in_external_connection.export
		input  wire        clk_clk,                                    //                                 clk.clk
		input  wire [3:0]  key_external_connection_export,             //             key_external_connection.export
		output wire        lcd_external_connection_RS,                 //             lcd_external_connection.RS
		output wire        lcd_external_connection_RW,                 //                                    .RW
		inout  wire [7:0]  lcd_external_connection_data,               //                                    .data
		output wire        lcd_external_connection_E,                  //                                    .E
		output wire [8:0]  ledg_external_connection_export,            //            ledg_external_connection.export
		output wire [17:0] ledr_external_connection_export,            //            ledr_external_connection.export
		input  wire        reset_reset_n,                              //                               reset.reset_n
		output wire [7:0]  sevseg_0_external_connection_export,        //        sevseg_0_external_connection.export
		output wire [7:0]  sevseg_1_external_connection_export,        //        sevseg_1_external_connection.export
		output wire [15:0] sevseg_2_external_connection_export,        //        sevseg_2_external_connection.export
		input  wire [9:0]  sw_external_connection_export               //              sw_external_connection.export
	);

	wire         nios2_qsys_debug_reset_request_reset;                      // nios2_qsys:debug_reset_request -> [camera_blue_in:reset_n, camera_green_in:reset_n, camera_red_in:reset_n, key:reset_n, lcd_0:reset_n, ledg:reset_n, ledr:reset_n, mm_interconnect_0:sysid_qsys_reset_reset_bridge_in_reset_reset, rst_controller:reset_in1, sevseg_0:reset_n, sevseg_1:reset_n, sevseg_2:reset_n, sw:reset_n, sysid_qsys:reset_n, timer:reset_n]
	wire  [31:0] nios2_qsys_data_master_readdata;                           // mm_interconnect_0:nios2_qsys_data_master_readdata -> nios2_qsys:d_readdata
	wire         nios2_qsys_data_master_waitrequest;                        // mm_interconnect_0:nios2_qsys_data_master_waitrequest -> nios2_qsys:d_waitrequest
	wire         nios2_qsys_data_master_debugaccess;                        // nios2_qsys:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_data_master_debugaccess
	wire  [19:0] nios2_qsys_data_master_address;                            // nios2_qsys:d_address -> mm_interconnect_0:nios2_qsys_data_master_address
	wire   [3:0] nios2_qsys_data_master_byteenable;                         // nios2_qsys:d_byteenable -> mm_interconnect_0:nios2_qsys_data_master_byteenable
	wire         nios2_qsys_data_master_read;                               // nios2_qsys:d_read -> mm_interconnect_0:nios2_qsys_data_master_read
	wire         nios2_qsys_data_master_write;                              // nios2_qsys:d_write -> mm_interconnect_0:nios2_qsys_data_master_write
	wire  [31:0] nios2_qsys_data_master_writedata;                          // nios2_qsys:d_writedata -> mm_interconnect_0:nios2_qsys_data_master_writedata
	wire  [31:0] nios2_qsys_instruction_master_readdata;                    // mm_interconnect_0:nios2_qsys_instruction_master_readdata -> nios2_qsys:i_readdata
	wire         nios2_qsys_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_qsys_instruction_master_waitrequest -> nios2_qsys:i_waitrequest
	wire  [18:0] nios2_qsys_instruction_master_address;                     // nios2_qsys:i_address -> mm_interconnect_0:nios2_qsys_instruction_master_address
	wire         nios2_qsys_instruction_master_read;                        // nios2_qsys:i_read -> mm_interconnect_0:nios2_qsys_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_control_slave_readdata;       // sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_control_slave_address;        // mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire   [7:0] mm_interconnect_0_lcd_0_control_slave_readdata;            // lcd_0:readdata -> mm_interconnect_0:lcd_0_control_slave_readdata
	wire   [1:0] mm_interconnect_0_lcd_0_control_slave_address;             // mm_interconnect_0:lcd_0_control_slave_address -> lcd_0:address
	wire         mm_interconnect_0_lcd_0_control_slave_read;                // mm_interconnect_0:lcd_0_control_slave_read -> lcd_0:read
	wire         mm_interconnect_0_lcd_0_control_slave_begintransfer;       // mm_interconnect_0:lcd_0_control_slave_begintransfer -> lcd_0:begintransfer
	wire         mm_interconnect_0_lcd_0_control_slave_write;               // mm_interconnect_0:lcd_0_control_slave_write -> lcd_0:write
	wire   [7:0] mm_interconnect_0_lcd_0_control_slave_writedata;           // mm_interconnect_0:lcd_0_control_slave_writedata -> lcd_0:writedata
	wire  [31:0] mm_interconnect_0_nios2_qsys_debug_mem_slave_readdata;     // nios2_qsys:debug_mem_slave_readdata -> mm_interconnect_0:nios2_qsys_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_qsys_debug_mem_slave_waitrequest;  // nios2_qsys:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_qsys_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_qsys_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_qsys_debug_mem_slave_debugaccess -> nios2_qsys:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_qsys_debug_mem_slave_address;      // mm_interconnect_0:nios2_qsys_debug_mem_slave_address -> nios2_qsys:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_qsys_debug_mem_slave_read;         // mm_interconnect_0:nios2_qsys_debug_mem_slave_read -> nios2_qsys:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_qsys_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_qsys_debug_mem_slave_byteenable -> nios2_qsys:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_qsys_debug_mem_slave_write;        // mm_interconnect_0:nios2_qsys_debug_mem_slave_write -> nios2_qsys:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_qsys_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_qsys_debug_mem_slave_writedata -> nios2_qsys:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_s1_chipselect;            // mm_interconnect_0:onchip_memory2_s1_chipselect -> onchip_memory2:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_readdata;              // onchip_memory2:readdata -> mm_interconnect_0:onchip_memory2_s1_readdata
	wire  [14:0] mm_interconnect_0_onchip_memory2_s1_address;               // mm_interconnect_0:onchip_memory2_s1_address -> onchip_memory2:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_s1_byteenable;            // mm_interconnect_0:onchip_memory2_s1_byteenable -> onchip_memory2:byteenable
	wire         mm_interconnect_0_onchip_memory2_s1_write;                 // mm_interconnect_0:onchip_memory2_s1_write -> onchip_memory2:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_writedata;             // mm_interconnect_0:onchip_memory2_s1_writedata -> onchip_memory2:writedata
	wire         mm_interconnect_0_onchip_memory2_s1_clken;                 // mm_interconnect_0:onchip_memory2_s1_clken -> onchip_memory2:clken
	wire         mm_interconnect_0_ledg_s1_chipselect;                      // mm_interconnect_0:ledg_s1_chipselect -> ledg:chipselect
	wire  [31:0] mm_interconnect_0_ledg_s1_readdata;                        // ledg:readdata -> mm_interconnect_0:ledg_s1_readdata
	wire   [1:0] mm_interconnect_0_ledg_s1_address;                         // mm_interconnect_0:ledg_s1_address -> ledg:address
	wire         mm_interconnect_0_ledg_s1_write;                           // mm_interconnect_0:ledg_s1_write -> ledg:write_n
	wire  [31:0] mm_interconnect_0_ledg_s1_writedata;                       // mm_interconnect_0:ledg_s1_writedata -> ledg:writedata
	wire  [31:0] mm_interconnect_0_sw_s1_readdata;                          // sw:readdata -> mm_interconnect_0:sw_s1_readdata
	wire   [1:0] mm_interconnect_0_sw_s1_address;                           // mm_interconnect_0:sw_s1_address -> sw:address
	wire  [31:0] mm_interconnect_0_key_s1_readdata;                         // key:readdata -> mm_interconnect_0:key_s1_readdata
	wire   [1:0] mm_interconnect_0_key_s1_address;                          // mm_interconnect_0:key_s1_address -> key:address
	wire         mm_interconnect_0_timer_s1_chipselect;                     // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                       // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                        // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                          // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                      // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire         mm_interconnect_0_sevseg_0_s1_chipselect;                  // mm_interconnect_0:sevseg_0_s1_chipselect -> sevseg_0:chipselect
	wire  [31:0] mm_interconnect_0_sevseg_0_s1_readdata;                    // sevseg_0:readdata -> mm_interconnect_0:sevseg_0_s1_readdata
	wire   [1:0] mm_interconnect_0_sevseg_0_s1_address;                     // mm_interconnect_0:sevseg_0_s1_address -> sevseg_0:address
	wire         mm_interconnect_0_sevseg_0_s1_write;                       // mm_interconnect_0:sevseg_0_s1_write -> sevseg_0:write_n
	wire  [31:0] mm_interconnect_0_sevseg_0_s1_writedata;                   // mm_interconnect_0:sevseg_0_s1_writedata -> sevseg_0:writedata
	wire         mm_interconnect_0_sevseg_1_s1_chipselect;                  // mm_interconnect_0:sevseg_1_s1_chipselect -> sevseg_1:chipselect
	wire  [31:0] mm_interconnect_0_sevseg_1_s1_readdata;                    // sevseg_1:readdata -> mm_interconnect_0:sevseg_1_s1_readdata
	wire   [1:0] mm_interconnect_0_sevseg_1_s1_address;                     // mm_interconnect_0:sevseg_1_s1_address -> sevseg_1:address
	wire         mm_interconnect_0_sevseg_1_s1_write;                       // mm_interconnect_0:sevseg_1_s1_write -> sevseg_1:write_n
	wire  [31:0] mm_interconnect_0_sevseg_1_s1_writedata;                   // mm_interconnect_0:sevseg_1_s1_writedata -> sevseg_1:writedata
	wire         mm_interconnect_0_sevseg_2_s1_chipselect;                  // mm_interconnect_0:sevseg_2_s1_chipselect -> sevseg_2:chipselect
	wire  [31:0] mm_interconnect_0_sevseg_2_s1_readdata;                    // sevseg_2:readdata -> mm_interconnect_0:sevseg_2_s1_readdata
	wire   [1:0] mm_interconnect_0_sevseg_2_s1_address;                     // mm_interconnect_0:sevseg_2_s1_address -> sevseg_2:address
	wire         mm_interconnect_0_sevseg_2_s1_write;                       // mm_interconnect_0:sevseg_2_s1_write -> sevseg_2:write_n
	wire  [31:0] mm_interconnect_0_sevseg_2_s1_writedata;                   // mm_interconnect_0:sevseg_2_s1_writedata -> sevseg_2:writedata
	wire         mm_interconnect_0_ledr_s1_chipselect;                      // mm_interconnect_0:ledr_s1_chipselect -> ledr:chipselect
	wire  [31:0] mm_interconnect_0_ledr_s1_readdata;                        // ledr:readdata -> mm_interconnect_0:ledr_s1_readdata
	wire   [1:0] mm_interconnect_0_ledr_s1_address;                         // mm_interconnect_0:ledr_s1_address -> ledr:address
	wire         mm_interconnect_0_ledr_s1_write;                           // mm_interconnect_0:ledr_s1_write -> ledr:write_n
	wire  [31:0] mm_interconnect_0_ledr_s1_writedata;                       // mm_interconnect_0:ledr_s1_writedata -> ledr:writedata
	wire  [31:0] mm_interconnect_0_camera_red_in_s1_readdata;               // camera_red_in:readdata -> mm_interconnect_0:camera_red_in_s1_readdata
	wire   [1:0] mm_interconnect_0_camera_red_in_s1_address;                // mm_interconnect_0:camera_red_in_s1_address -> camera_red_in:address
	wire  [31:0] mm_interconnect_0_camera_green_in_s1_readdata;             // camera_green_in:readdata -> mm_interconnect_0:camera_green_in_s1_readdata
	wire   [1:0] mm_interconnect_0_camera_green_in_s1_address;              // mm_interconnect_0:camera_green_in_s1_address -> camera_green_in:address
	wire  [31:0] mm_interconnect_0_camera_blue_in_s1_readdata;              // camera_blue_in:readdata -> mm_interconnect_0:camera_blue_in_s1_readdata
	wire   [1:0] mm_interconnect_0_camera_blue_in_s1_address;               // mm_interconnect_0:camera_blue_in_s1_address -> camera_blue_in:address
	wire         irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // timer:irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_qsys_irq_irq;                                        // irq_mapper:sender_irq -> nios2_qsys:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:nios2_qsys_reset_reset_bridge_in_reset_reset, nios2_qsys:reset_n, onchip_memory2:reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [nios2_qsys:reset_req, onchip_memory2:reset_req, rst_translator:reset_req_in]

	DE2_115_QSYS_camera_blue_in camera_blue_in (
		.clk      (clk_clk),                                      //                 clk.clk
		.reset_n  (~nios2_qsys_debug_reset_request_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_camera_blue_in_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_camera_blue_in_s1_readdata), //                    .readdata
		.in_port  (camera_blue_in_external_connection_export)     // external_connection.export
	);

	DE2_115_QSYS_camera_blue_in camera_green_in (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~nios2_qsys_debug_reset_request_reset),         //               reset.reset_n
		.address  (mm_interconnect_0_camera_green_in_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_camera_green_in_s1_readdata), //                    .readdata
		.in_port  (camera_green_in_external_connection_export)     // external_connection.export
	);

	DE2_115_QSYS_camera_blue_in camera_red_in (
		.clk      (clk_clk),                                     //                 clk.clk
		.reset_n  (~nios2_qsys_debug_reset_request_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_camera_red_in_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_camera_red_in_s1_readdata), //                    .readdata
		.in_port  (camera_red_in_external_connection_export)     // external_connection.export
	);

	DE2_115_QSYS_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	DE2_115_QSYS_key key (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~nios2_qsys_debug_reset_request_reset), //               reset.reset_n
		.address  (mm_interconnect_0_key_s1_address),      //                  s1.address
		.readdata (mm_interconnect_0_key_s1_readdata),     //                    .readdata
		.in_port  (key_external_connection_export)         // external_connection.export
	);

	DE2_115_QSYS_lcd_0 lcd_0 (
		.reset_n       (~nios2_qsys_debug_reset_request_reset),               //         reset.reset_n
		.clk           (clk_clk),                                             //           clk.clk
		.begintransfer (mm_interconnect_0_lcd_0_control_slave_begintransfer), // control_slave.begintransfer
		.read          (mm_interconnect_0_lcd_0_control_slave_read),          //              .read
		.write         (mm_interconnect_0_lcd_0_control_slave_write),         //              .write
		.readdata      (mm_interconnect_0_lcd_0_control_slave_readdata),      //              .readdata
		.writedata     (mm_interconnect_0_lcd_0_control_slave_writedata),     //              .writedata
		.address       (mm_interconnect_0_lcd_0_control_slave_address),       //              .address
		.LCD_RS        (lcd_external_connection_RS),                          //      external.export
		.LCD_RW        (lcd_external_connection_RW),                          //              .export
		.LCD_data      (lcd_external_connection_data),                        //              .export
		.LCD_E         (lcd_external_connection_E)                            //              .export
	);

	DE2_115_QSYS_ledg ledg (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~nios2_qsys_debug_reset_request_reset), //               reset.reset_n
		.address    (mm_interconnect_0_ledg_s1_address),     //                  s1.address
		.write_n    (~mm_interconnect_0_ledg_s1_write),      //                    .write_n
		.writedata  (mm_interconnect_0_ledg_s1_writedata),   //                    .writedata
		.chipselect (mm_interconnect_0_ledg_s1_chipselect),  //                    .chipselect
		.readdata   (mm_interconnect_0_ledg_s1_readdata),    //                    .readdata
		.out_port   (ledg_external_connection_export)        // external_connection.export
	);

	DE2_115_QSYS_ledr ledr (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~nios2_qsys_debug_reset_request_reset), //               reset.reset_n
		.address    (mm_interconnect_0_ledr_s1_address),     //                  s1.address
		.write_n    (~mm_interconnect_0_ledr_s1_write),      //                    .write_n
		.writedata  (mm_interconnect_0_ledr_s1_writedata),   //                    .writedata
		.chipselect (mm_interconnect_0_ledr_s1_chipselect),  //                    .chipselect
		.readdata   (mm_interconnect_0_ledr_s1_readdata),    //                    .readdata
		.out_port   (ledr_external_connection_export)        // external_connection.export
	);

	DE2_115_QSYS_nios2_qsys nios2_qsys (
		.clk                                 (clk_clk),                                                  //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                          //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                       //                          .reset_req
		.d_address                           (nios2_qsys_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_qsys_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_qsys_data_master_read),                              //                          .read
		.d_readdata                          (nios2_qsys_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_qsys_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_qsys_data_master_write),                             //                          .write
		.d_writedata                         (nios2_qsys_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_qsys_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_qsys_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_qsys_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_qsys_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_qsys_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_qsys_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_qsys_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_qsys_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_qsys_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_qsys_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_qsys_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_qsys_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_qsys_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_qsys_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_qsys_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                          // custom_instruction_master.readra
	);

	DE2_115_QSYS_onchip_memory2 onchip_memory2 (
		.clk        (clk_clk),                                        //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                 // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),             //       .reset_req
		.freeze     (1'b0)                                            // (terminated)
	);

	DE2_115_QSYS_sevseg_0 sevseg_0 (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~nios2_qsys_debug_reset_request_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_sevseg_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sevseg_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sevseg_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sevseg_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sevseg_0_s1_readdata),   //                    .readdata
		.out_port   (sevseg_0_external_connection_export)       // external_connection.export
	);

	DE2_115_QSYS_sevseg_0 sevseg_1 (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~nios2_qsys_debug_reset_request_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_sevseg_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sevseg_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sevseg_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sevseg_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sevseg_1_s1_readdata),   //                    .readdata
		.out_port   (sevseg_1_external_connection_export)       // external_connection.export
	);

	DE2_115_QSYS_sevseg_2 sevseg_2 (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~nios2_qsys_debug_reset_request_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_sevseg_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sevseg_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sevseg_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sevseg_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sevseg_2_s1_readdata),   //                    .readdata
		.out_port   (sevseg_2_external_connection_export)       // external_connection.export
	);

	DE2_115_QSYS_sw sw (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~nios2_qsys_debug_reset_request_reset), //               reset.reset_n
		.address  (mm_interconnect_0_sw_s1_address),       //                  s1.address
		.readdata (mm_interconnect_0_sw_s1_readdata),      //                    .readdata
		.in_port  (sw_external_connection_export)          // external_connection.export
	);

	DE2_115_QSYS_sysid_qsys sysid_qsys (
		.clock    (clk_clk),                                             //           clk.clk
		.reset_n  (~nios2_qsys_debug_reset_request_reset),               //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_control_slave_address)   //              .address
	);

	DE2_115_QSYS_timer timer (
		.clk        (clk_clk),                               //   clk.clk
		.reset_n    (~nios2_qsys_debug_reset_request_reset), // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)               //   irq.irq
	);

	DE2_115_QSYS_mm_interconnect_0 mm_interconnect_0 (
		.clk_50_clk_clk                               (clk_clk),                                                   //                             clk_50_clk.clk
		.nios2_qsys_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // nios2_qsys_reset_reset_bridge_in_reset.reset
		.sysid_qsys_reset_reset_bridge_in_reset_reset (nios2_qsys_debug_reset_request_reset),                      // sysid_qsys_reset_reset_bridge_in_reset.reset
		.nios2_qsys_data_master_address               (nios2_qsys_data_master_address),                            //                 nios2_qsys_data_master.address
		.nios2_qsys_data_master_waitrequest           (nios2_qsys_data_master_waitrequest),                        //                                       .waitrequest
		.nios2_qsys_data_master_byteenable            (nios2_qsys_data_master_byteenable),                         //                                       .byteenable
		.nios2_qsys_data_master_read                  (nios2_qsys_data_master_read),                               //                                       .read
		.nios2_qsys_data_master_readdata              (nios2_qsys_data_master_readdata),                           //                                       .readdata
		.nios2_qsys_data_master_write                 (nios2_qsys_data_master_write),                              //                                       .write
		.nios2_qsys_data_master_writedata             (nios2_qsys_data_master_writedata),                          //                                       .writedata
		.nios2_qsys_data_master_debugaccess           (nios2_qsys_data_master_debugaccess),                        //                                       .debugaccess
		.nios2_qsys_instruction_master_address        (nios2_qsys_instruction_master_address),                     //          nios2_qsys_instruction_master.address
		.nios2_qsys_instruction_master_waitrequest    (nios2_qsys_instruction_master_waitrequest),                 //                                       .waitrequest
		.nios2_qsys_instruction_master_read           (nios2_qsys_instruction_master_read),                        //                                       .read
		.nios2_qsys_instruction_master_readdata       (nios2_qsys_instruction_master_readdata),                    //                                       .readdata
		.camera_blue_in_s1_address                    (mm_interconnect_0_camera_blue_in_s1_address),               //                      camera_blue_in_s1.address
		.camera_blue_in_s1_readdata                   (mm_interconnect_0_camera_blue_in_s1_readdata),              //                                       .readdata
		.camera_green_in_s1_address                   (mm_interconnect_0_camera_green_in_s1_address),              //                     camera_green_in_s1.address
		.camera_green_in_s1_readdata                  (mm_interconnect_0_camera_green_in_s1_readdata),             //                                       .readdata
		.camera_red_in_s1_address                     (mm_interconnect_0_camera_red_in_s1_address),                //                       camera_red_in_s1.address
		.camera_red_in_s1_readdata                    (mm_interconnect_0_camera_red_in_s1_readdata),               //                                       .readdata
		.jtag_uart_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //            jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                       .write
		.jtag_uart_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                       .read
		.jtag_uart_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                       .readdata
		.jtag_uart_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                       .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                       .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                       .chipselect
		.key_s1_address                               (mm_interconnect_0_key_s1_address),                          //                                 key_s1.address
		.key_s1_readdata                              (mm_interconnect_0_key_s1_readdata),                         //                                       .readdata
		.lcd_0_control_slave_address                  (mm_interconnect_0_lcd_0_control_slave_address),             //                    lcd_0_control_slave.address
		.lcd_0_control_slave_write                    (mm_interconnect_0_lcd_0_control_slave_write),               //                                       .write
		.lcd_0_control_slave_read                     (mm_interconnect_0_lcd_0_control_slave_read),                //                                       .read
		.lcd_0_control_slave_readdata                 (mm_interconnect_0_lcd_0_control_slave_readdata),            //                                       .readdata
		.lcd_0_control_slave_writedata                (mm_interconnect_0_lcd_0_control_slave_writedata),           //                                       .writedata
		.lcd_0_control_slave_begintransfer            (mm_interconnect_0_lcd_0_control_slave_begintransfer),       //                                       .begintransfer
		.ledg_s1_address                              (mm_interconnect_0_ledg_s1_address),                         //                                ledg_s1.address
		.ledg_s1_write                                (mm_interconnect_0_ledg_s1_write),                           //                                       .write
		.ledg_s1_readdata                             (mm_interconnect_0_ledg_s1_readdata),                        //                                       .readdata
		.ledg_s1_writedata                            (mm_interconnect_0_ledg_s1_writedata),                       //                                       .writedata
		.ledg_s1_chipselect                           (mm_interconnect_0_ledg_s1_chipselect),                      //                                       .chipselect
		.ledr_s1_address                              (mm_interconnect_0_ledr_s1_address),                         //                                ledr_s1.address
		.ledr_s1_write                                (mm_interconnect_0_ledr_s1_write),                           //                                       .write
		.ledr_s1_readdata                             (mm_interconnect_0_ledr_s1_readdata),                        //                                       .readdata
		.ledr_s1_writedata                            (mm_interconnect_0_ledr_s1_writedata),                       //                                       .writedata
		.ledr_s1_chipselect                           (mm_interconnect_0_ledr_s1_chipselect),                      //                                       .chipselect
		.nios2_qsys_debug_mem_slave_address           (mm_interconnect_0_nios2_qsys_debug_mem_slave_address),      //             nios2_qsys_debug_mem_slave.address
		.nios2_qsys_debug_mem_slave_write             (mm_interconnect_0_nios2_qsys_debug_mem_slave_write),        //                                       .write
		.nios2_qsys_debug_mem_slave_read              (mm_interconnect_0_nios2_qsys_debug_mem_slave_read),         //                                       .read
		.nios2_qsys_debug_mem_slave_readdata          (mm_interconnect_0_nios2_qsys_debug_mem_slave_readdata),     //                                       .readdata
		.nios2_qsys_debug_mem_slave_writedata         (mm_interconnect_0_nios2_qsys_debug_mem_slave_writedata),    //                                       .writedata
		.nios2_qsys_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_qsys_debug_mem_slave_byteenable),   //                                       .byteenable
		.nios2_qsys_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_qsys_debug_mem_slave_waitrequest),  //                                       .waitrequest
		.nios2_qsys_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_qsys_debug_mem_slave_debugaccess),  //                                       .debugaccess
		.onchip_memory2_s1_address                    (mm_interconnect_0_onchip_memory2_s1_address),               //                      onchip_memory2_s1.address
		.onchip_memory2_s1_write                      (mm_interconnect_0_onchip_memory2_s1_write),                 //                                       .write
		.onchip_memory2_s1_readdata                   (mm_interconnect_0_onchip_memory2_s1_readdata),              //                                       .readdata
		.onchip_memory2_s1_writedata                  (mm_interconnect_0_onchip_memory2_s1_writedata),             //                                       .writedata
		.onchip_memory2_s1_byteenable                 (mm_interconnect_0_onchip_memory2_s1_byteenable),            //                                       .byteenable
		.onchip_memory2_s1_chipselect                 (mm_interconnect_0_onchip_memory2_s1_chipselect),            //                                       .chipselect
		.onchip_memory2_s1_clken                      (mm_interconnect_0_onchip_memory2_s1_clken),                 //                                       .clken
		.sevseg_0_s1_address                          (mm_interconnect_0_sevseg_0_s1_address),                     //                            sevseg_0_s1.address
		.sevseg_0_s1_write                            (mm_interconnect_0_sevseg_0_s1_write),                       //                                       .write
		.sevseg_0_s1_readdata                         (mm_interconnect_0_sevseg_0_s1_readdata),                    //                                       .readdata
		.sevseg_0_s1_writedata                        (mm_interconnect_0_sevseg_0_s1_writedata),                   //                                       .writedata
		.sevseg_0_s1_chipselect                       (mm_interconnect_0_sevseg_0_s1_chipselect),                  //                                       .chipselect
		.sevseg_1_s1_address                          (mm_interconnect_0_sevseg_1_s1_address),                     //                            sevseg_1_s1.address
		.sevseg_1_s1_write                            (mm_interconnect_0_sevseg_1_s1_write),                       //                                       .write
		.sevseg_1_s1_readdata                         (mm_interconnect_0_sevseg_1_s1_readdata),                    //                                       .readdata
		.sevseg_1_s1_writedata                        (mm_interconnect_0_sevseg_1_s1_writedata),                   //                                       .writedata
		.sevseg_1_s1_chipselect                       (mm_interconnect_0_sevseg_1_s1_chipselect),                  //                                       .chipselect
		.sevseg_2_s1_address                          (mm_interconnect_0_sevseg_2_s1_address),                     //                            sevseg_2_s1.address
		.sevseg_2_s1_write                            (mm_interconnect_0_sevseg_2_s1_write),                       //                                       .write
		.sevseg_2_s1_readdata                         (mm_interconnect_0_sevseg_2_s1_readdata),                    //                                       .readdata
		.sevseg_2_s1_writedata                        (mm_interconnect_0_sevseg_2_s1_writedata),                   //                                       .writedata
		.sevseg_2_s1_chipselect                       (mm_interconnect_0_sevseg_2_s1_chipselect),                  //                                       .chipselect
		.sw_s1_address                                (mm_interconnect_0_sw_s1_address),                           //                                  sw_s1.address
		.sw_s1_readdata                               (mm_interconnect_0_sw_s1_readdata),                          //                                       .readdata
		.sysid_qsys_control_slave_address             (mm_interconnect_0_sysid_qsys_control_slave_address),        //               sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata            (mm_interconnect_0_sysid_qsys_control_slave_readdata),       //                                       .readdata
		.timer_s1_address                             (mm_interconnect_0_timer_s1_address),                        //                               timer_s1.address
		.timer_s1_write                               (mm_interconnect_0_timer_s1_write),                          //                                       .write
		.timer_s1_readdata                            (mm_interconnect_0_timer_s1_readdata),                       //                                       .readdata
		.timer_s1_writedata                           (mm_interconnect_0_timer_s1_writedata),                      //                                       .writedata
		.timer_s1_chipselect                          (mm_interconnect_0_timer_s1_chipselect)                      //                                       .chipselect
	);

	DE2_115_QSYS_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios2_qsys_irq_irq)              //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                       // reset_in0.reset
		.reset_in1      (nios2_qsys_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                              //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),       // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),   //          .reset_req
		.reset_req_in0  (1'b0),                                 // (terminated)
		.reset_req_in1  (1'b0),                                 // (terminated)
		.reset_in2      (1'b0),                                 // (terminated)
		.reset_req_in2  (1'b0),                                 // (terminated)
		.reset_in3      (1'b0),                                 // (terminated)
		.reset_req_in3  (1'b0),                                 // (terminated)
		.reset_in4      (1'b0),                                 // (terminated)
		.reset_req_in4  (1'b0),                                 // (terminated)
		.reset_in5      (1'b0),                                 // (terminated)
		.reset_req_in5  (1'b0),                                 // (terminated)
		.reset_in6      (1'b0),                                 // (terminated)
		.reset_req_in6  (1'b0),                                 // (terminated)
		.reset_in7      (1'b0),                                 // (terminated)
		.reset_req_in7  (1'b0),                                 // (terminated)
		.reset_in8      (1'b0),                                 // (terminated)
		.reset_req_in8  (1'b0),                                 // (terminated)
		.reset_in9      (1'b0),                                 // (terminated)
		.reset_req_in9  (1'b0),                                 // (terminated)
		.reset_in10     (1'b0),                                 // (terminated)
		.reset_req_in10 (1'b0),                                 // (terminated)
		.reset_in11     (1'b0),                                 // (terminated)
		.reset_req_in11 (1'b0),                                 // (terminated)
		.reset_in12     (1'b0),                                 // (terminated)
		.reset_req_in12 (1'b0),                                 // (terminated)
		.reset_in13     (1'b0),                                 // (terminated)
		.reset_req_in13 (1'b0),                                 // (terminated)
		.reset_in14     (1'b0),                                 // (terminated)
		.reset_req_in14 (1'b0),                                 // (terminated)
		.reset_in15     (1'b0),                                 // (terminated)
		.reset_req_in15 (1'b0)                                  // (terminated)
	);

endmodule
