��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���麍�Ks�%$����+d7��/��������ߔ,���<�E�]��&��z>��>�X�����`��B�㓪F:��ew���@�C�k�.U6�vά1�xrl9��Sr?$R�t��M��~3pwd��<�i��w_�)4ޟo$#)����4F�1s[�p;��Q�!��x44S�"s
S������D^q_\�e�k`�R<��H8��{Y�~|@�d�SGbUP��Ζ^\�w�QIx=�R�x���.�"����.��|4�z��.a'h�!��j0�ՙ ��M�q��3/V0Z>.�r�;;t���6�G����r�����,ڗ�#w�~�}	:��7˽|�}�+o��s?|�1#&���ֵ��EN�w���YF5��o��	y���m9E;��\u=�M���6H ��ђ2ט0�)�-����7�*gyb ݄Z:z<7���/��;�R����m�Ӏ ����ouY u<W�h���ȑ�n�� l-��cgN05{�PM��"�$C�oZaQ��ܤ:ͥ\��}�A�8HZ��¢-�Db(D�N��xQ\X�`�{�Z[b#C�0ڌhS��SV<�l��V%���e����G�$�̍�m����K`H�4=�Z�W(�.�5�db�-V���Y���z��^=�]l��X�rCJ*����&`:Z��#{ۄ"<��_~�e;�W�-&u��YKH�p�,Y��'�̞��c��j[(8�}���m���\5��g,/�$���� ��?���i�sE�f�J�w�����^K~]y\_��e,a�pB(�U�1U�Ol�4���b�OY�j�/�I)٣m�B��L��Ѓ���?+ʹ$TLnD�C�'�������2�T�O�ؐ���!����N9dм*��?�L�J��M��PԐQj��s�u���%*�'��Z΀B������d�E[��d ��LͿ��ǿ�	�~M�~������P�սWR��
�B���^��˦L����~�&z�~�{Ě� ���T�$������z>ӂ�`��8S[4�˔mh�nԯ��sm(C�Z��*\���߄�%.���G�S�}V����j�U�v	��,�{2��4�T� ^�@�����I��KUtL���Eˣf��~l��6dVJ)_�Uʎu?�2�btRfV�mlې�I�(>���?�,e����enŁ�."��ƅ���F���a�W��0ay�Y[��U�'=N��H �q��MT5�I�L�Fᬩ?F��:�ah\��;�~g�ϒ��+�.6�����s�Ϝ�hL�R]k�Y�B��N3KWU��'z[6����SCL/�Ԗ��??
�X��-}��a`��2�E���j��FQ����,cvk	�,��Y)�	c1��鐭��aa�sx�ƻ�w���̿�d�m݊p?}�$��_��/~��q:�}qc�Oyq��"��@+�+E�����}H��}�m�6(��{���|hQ`�����z[q�-�#�U�"<�&�������� ��e�?��eb)�⛙��s~�9����.�e���* ƿ��N�3^-�?�n��܀��m(�G�^�Z��*E�.�g��j��!�GQg�K���r��?*���$<8�H��%�i�,9�_�:3v�|ļۑ���|H�{v�t�}	oG�������;꫸�Y���7��:[���0�.90��5�������������B����O>;�Ģ0B�|�imڇpP`Q���](�2����uQj}�s�$"���~"����ǛpL�����$�j�b�"�J� �[3"�c������{�I�PڙPKa(�� K�P�t�kk.��V�hήi,�jϭ����z�$X�,&���ͲX���{14/-�b3�f���Dk�|g��K5�Aъ%���A�a^�%Z%�xʜ%z��zV]�}0�Զd�\q	�U����[���K��&gQ��
��M��$7>R��O!?�B:[�p�^=��hWf��COj�)���Rҳ$���_��tO��$��Ӝ ��D-�T��_�)�d�����ꩰ��5I@k�d[��0 :����a�_9��H�-�M�?���>��D$���F����Q��̶����x:9�#��ưR��UZ)���<z�b���x�Z�9dyT~�����o		�2�ԍ���~�r���^y�R!��EL�sJ)ޙ�ׁt��4~����Љ�/��T�'�χeŜWvM�g�����"CP���vTZ�)�����,��
�w$���дyP\��JJE��x��QDM׵oq+�k���鼣"پʇ0�ڗ¯��zY����i;ф��)g��[���r^�u�r�{&d>�����]�S7y������ێ����-�Aّ	;6u�a��(�VX�n��ɬQ�� g�Sf|@V�Xe�w����rߕ�� w������C���~����r�\�x��`P��U�ʱ2�쫰�ɏ�fÑ�
r�Ņ�}^�K�o(�@���M��G;�E	��;#��4��c����F9TX�d� eJ�(�XV��Sm�(�Yl��VB�s�|��-��JT�
�:�yk��R����w8mPE����&��v���i�;�/u��/�ê�-p;�
BJ��Y�)�_�q���_�s�{r�IؒT�ćh��K���!v'W+nQ�Sc���i�ĥx�`��o�LNXEmʦ�^�W�{_+"z����Ĩ����}2�W��|����J����Mz/��z>�>.��TR7����9��(�
�G�e��ņnԆ��DЛ{��-��?���p4ck9�1K]c"��
%3Q;��"b�u;N�۝��=B8ך~mNQ�y�G?�qP�#9��G!���ܩ*n��&-������jTS�D5�(�]�m����ɶx�����0�i-c�Z�wȓ
�x��E�#�������98;�|-汭G�����1����dC�,]WT�M�.�D��e��H�fo��2����!�gw�}��ߘ���q��9��ԘwĜ�ן�z>���v�$y}��`�%�ϖ��ZX�%�E��]��9H��p׎L�+�`�� ����=6�;jQ�Иa)�PN:㯼�����Gn>�,$S��b?�N]�
�G�J�h�L�yڔz�o��`��W��R���N9=���~=�,�k��d%����P�!�Foc��0Q4��h���],+�ٽ:}ٯ��G M�b*���w���c��Z�[9�ۋ�kJ��ʣ%5�i��X#�X���
���L�S'GVz���$P�5��a�v����y;2�.�K|S�B��ߟ5�Z�]?%����ƣZۙ.$�Ey�z��>����~��1C��`N�Q�l^g��q���n�����#������Arz�Ev<Y������<�ˀ�O�ПݮI�"��7�I*�`t�����s.�[������8�	�c2F�YNQ�1P��\7�j��/J�Dѣ�~M�{�$K9��#��D!-I�%ܺ�@����V�		\D(ͬMoItWD��oM:lm����wLs��͂�M�V��r���N��gh��o�C8,�3�n@����A��tϪ.�b�#�P7�L=*�}iM�.8&���RAi�RYÏ#w��oy�R�$�X��dq�	H�߶lI��U/ȡ�KB�m�����z|�<�r'�M�H��UW*�F����` �o/���a�>.Y�u+��}:@�"�[0�	�WW�%I}>�@v��1�USE���ʿL�ٚ�6��aOv�	V���EHԥ)��H�؂�(밼�<b�L~X�?t0� M!���|iS��9��W`��o?�� ������k��%g>{5Ǧ�ɉBd�˚&S�vΩ3�Bp'�)P�����!�@��'���]�}}��N/��*H偒��镲�^�L3���Ůs-�]��������%�)}�Տ���:�y�	]�u"�s�L��榰B֛"��L�O����ϔ[��i4K�5-�jN!����rC(�X�64�Fv�E��&~��1�T�-į*W���Tu�F�>�C��xo��M�*��ؓ*+6����σ ����������.<�i�`��ս�L�N����bK�ƕüL��+�3�Y��]~��>�u�{&�V5�$d�i�v~�?Vtli�k}��_�mBłbi���H"����XL9`��7?j쨺C�:��;G�V�ɓ�5�Ff��w�n�LPc/����1J����^\��*��|_D+�93m�-�7�+���AM{���$O�eD���cd�j�~�ݿ;���*�|z�=.�JlfR�S������~Ma� ^��Ph�oJ&��k���C� ��]�������/�I��0����WhnX�"0D�`��<��*���,��P�n��Q�E�Y}?AGZ�� .;��b�h��I7� ה�DQ]��c�Q��Z.�n� U��\�m��M|-�� ����Oܐ��5aV�Q�S�C�pF}��<�=DS9XVڀ�sRN���2ύ�LgO�L$ uĐ���ԅh-��+�;zm{ś�P���{s����{ߟ4���س�Mh��6��5Oŉw�?F�����s�<󓩿�*VWOd.�$������bf]��"��LD�Tޫ>Ǧ�o��M|��̅� W~� �y@[�{�*��/"2g��������)c!����cJ�jY�����v[L��s��sT=B��>cR�
��y�f
���]�V=p�:Nh2�w��z��'�w:kpý0w9F.7Q\#-j�n��D�]/��B��H��\�((8^t)勪̠�ȁ����x82H�p+���=����㝜	��d���F�f�?ӡ�8�T���>T5��l٩G���f�7�!�e�,E2�Ȩ{�H_�p�<'�Y��t'�{3���L[>i-���ߤT����*�[<rJ*u��b"���/�),\��/{4�@�o�#:��}2�)��uU�TA�e��hu���y����4�)�	�4���ը��j�2�q�u#b����v ��D�8Й i��Tr���i�n�
1s��_��30�+�>�/O{�j��,�ujz�rqI��oWOv(K�,���3�j��,���jt"}4��3��e\*�\�9*ܔq�6�n0S/�����
�Uѱ�_��8����K�����'��	2&z?bV�^�E��@�F��O�U��P�;+�Y@E��>\��,GY_��n�7(%m.Z�|�L���(��h2�6�
��~W�9W_A����1�@!oVt���l�>�+kג�Oo�mJ!�Mq�>����S���«�0�>�!��f�o�"N�X��'z��Zq�gF.�>��2,_�c�V}�8�#]HM��� q������$�#lO��.����=R	�Ƌ���0�O�����?�;l0x��^��������`Y�c%K�I��T4PD4w�ƈ�@Vsn�n�D��!ף���QeP:�>��H��J�BL�yS� (����$T��A��{���F*q�m��{qQ��l��#�%?�j˂�^�!�a�����E��f�O1����T��a��~O�N���$�sC�0��8�D Q\~+CVS?������E��g��fL�Fl���Y��h�+%,	[:�dXY������O�lr<-�_��H�?�CosZ�d�G�-؀Mn�����������uXI~!a'���S1�����k`��z�9����x��h�E�mPIo�&q��<Ɍ?1D�I�H�@Mbu�q��,�aV�����e�p��;t�w�,V�Nڽ�k���;��0�d���n^F�9	�4a����k���,@���X���u�Bˉ�ں},���u�.8cU^�u��Х-9��E��q'0��Zk@�s��G��w�g9�X'e�oX]�A��*������ϗ�����~ʢ���_���9Z����q�1��%�
��K�EiW93��|Hv�0�ξW��
	0��X��1@���J����a��v���[тd7���(M� �r\�^���Qc�C$֢�)09�2�OT�H��y�K��#�R�鶂J�NMT��0��b|Ư��Zq���{��q#���O�;b�O)�y�aR��ZCw����WU`9��t����� 2K�,o���^����`2?�6N\�k]c�^L:4:xIֵ��Sژ.W��p2Q����+�t���(�VZ�&�?�ߋ{��	>�,�@�
�T�5�T�H�&j�E�O�d�ɛeeƄ�nՇ,��-��P�;{�`�5}P��k�ng�N�7@��3���
�]׃��~�ݧ����l��wT��X_���&bXQ��'�:�6�v��ߝ�(�D�]�.��,#�#�ȧ���a�d3�;�,Kp�թP$�E��n/gpsGen�ƣ�*}Ϡ��Z2��n�	R�+8
M\Z/�uv,�:%�����?�� ̄��}�D�w�����X�Q�2Xa��]��g���>���R5>ם�ݺa-�
8���W�� l��L��h
Ui���2ƃ�^�e�N����:��ay�xּ�cEkc.=���{�]�HG��ݝ�i�*�غ:�a��ow�ꫭ�L�F/��u�k�dK�� �9��g�.`��4��*�#�b���m��ڛuh������EMY����Z�~#g0�^xA�$�����g������/�s9U�fzN�ړ�jD���m�K�c����r��t����f�r�0#� �=����J̒����j���5�C�W��w�z4���Q�:i�b���m#�C���y`9�D�~�z�8��|j��!n���q��ˑ��X${�T�����f���E�@i]�*J_�^���>��Wu6I�]D͙s/"*�S�ram���nk\<��	��8��ϥ!z��:���Ϲz$�W���W�2����V��jQ?������˶�z�U�M�a#Po�}R��[�u2��ݛ����m�o���+.�d*6���p��\���d\z�01���\+����tZ����.)�q��أ`��#(�U�����WB������2��	�wO�+{f:�L�oy���t�g�s�$���^}��+����FiM,�Ԗ�ʞ�ج�5a-x�ۋ��aZ�E��kB��Ŏ*O�jDV������&bn�97���/,�6@,GHob,M7�!���J�;�G�F�dZ�.X�ѯ�N�0����,��e�i�93.M�̪���Of�8w�_8wR�����~*g��%����srm�a�>�iH��%����NsY�v�2�XD�?o��I�a0�M�.(��<>g��V��}�%"��M�0�2��@��fc���mq�Ӏ��m���$�}��?� �X�g�eVb���2k�EB~�qOb)���:O�}���u��e�����%���~!���H}eݵ��-�ﳜ�uF�/;d�Ȏ���2��dsHj�94�����PFx�ʹ�5$Ϭ�ISJ�`�+<����ƍj=�ۦG}��r�~��q��{�V�:���%"��_nzDG�*Xéé�nr�{q;Uy��F'i2(���fo�<o^��!�Yiز����FԶ6�G��Ċ57��w�h�q��;ڢ&�U��y�T��e B��j��94EGhZ�[i>�X�w������TEѯy�+�������,���Y�0 VA�\*���Vj?��l��rQ#��&�~qF9��`U�!�>ǥ+%9�)�z�K����e�N�w��{�.辒(NΎ;$��i�B�M�B�����Ad�]5�ҿ�g�	�]C�A����J�e���g�(�#��<����+��vr�]ΨKV��.�a��f���π�@��0=�=*5�E�GgMX���!�4�֍8o�CಳM���k_��u���5g:�����HC��y���o���D��r�v0���Q2�"��Ĵ5���A���Sv�c����F
Ԡ��L�g�z�Gx���`�Ԯ|��%f]{Gts�5�����I��e/c~�✌�B϶sE����5O��c��+�fY��noj�K�}�G�2�Mu�dcK�+��^���TF�sb1�I��9Wq�ns�W	�XJ0���X�A=�Ct0����+�eG����|ǎ�NO��$�0|��Ә��Fw�bY�l��t,��4�B���hWp:���.�T<}��p�R��2-�w"�O��+���ϕ�X2��E�|�r��O��� ��l.�4���Ǎ��Vz���iK�^Ӧ��1?Db����l��r_�"�+�hic�o�q��Zx�w:��q����?����ug$��x0�е���XYA���bp��$���zoa���,"^�Mqc�s�ͭD�7��o�͞ :���N�B��({�oy��]'31oO8�{�_&/+�zS{]V[Q�� A�K���/�xx|���ZF�\�x����t�r�%Z#�톺�-. ,x$Ҍ��6���N��b]%ށ���4�Nt�������>uW�2cn���2'�<a�	�XZ+���E�7T��
X����=�M���a6�.D��Go�9��� �<38.=B�	qyb��t�lm���aE�&bl�2�^D5W�%!���8�v��
+�{�jKm;���͏�a��A��6�F/P�>��a�2˼��r89�V6[S5�cl<+��?g�b��<�)
��u��.���pb�=D��8k�ev��|�L���I����L�m�
G�jK��o@P��x|��1�N1[Za/	d��F,�Pϡ����j�2����4X�Ǡ}/��Z�3FM��0,�eBu�C���<n\n�{M�F�9�ȢH��0�(��u9#�Բ�-M}m�p��X�v�vV���tlx��*�5k�/�j�n��;��9bٗ�@D��ړ�x?�5�9��U����v��?SIEǟ��*�L
��`vPX��VrsR�5RYC�b��I7@ZY�P���\�c��d,����N`�i�d�.����(��]:v'��|1�ڐ��S�!�9�~b��rMQ�w��x���)0��1f��%�5G�kQd�
{��I��9��b�
�UdH���F�0��p�l��?�t�̖`>���RkŅ�fd��FWB�)CKL&d-E�/�e��������E��fY���9YA��x#��g�R4w�
��ͮX����tǢEO�7��N�NK<P�5@F�����?/vĢ��X�WO� ��W��ە�!�����w��:+�Ͱ'p�Wrؿ�)��/�ʕ����n��v����gK���x�!�rJv���`�N����p>�s�A��O20�r��y9�o{�����%"FTį���|ȫ�Y; hM��y��=\4����i�699i`!�r�K�����!�����aT���SQ���ª��8��*^�����T/��;\6:u�J͂�C-Z�+/O\�#���F<��e +��2��p���$�G"���\�Ƙh��j��z#��8�!�1)����4�c�y<F �,��[/��}�(���ט�o����� \����^��e�OM�Z�4���p����m
��6Sو�DU�}���ܽh� �sH��h(��\M����|3���O���֛}V�q��x��]C�l���ŗy�{p���ӑ�t�t0
r��eA�~F=͠M��
6��A��+�ͳ8!w��Ȱ���E�S�m�y���w�������\T�5�UȅL���=/|�b#�����P[P_>`�����-��t�m�0��"�j�m!p8����]y����6��Xfo�M�Ǐ��8z�������Un�p��ø�o�l�dڼz��n"P�\���$�(a���W����'*O�t��{�6em�Q���]�d�:�L7#��-�Q�����k��*W��el��'D�w�^����k�\0�n�B���\�=v; |��,��l�ۍtD���:���ޙ��r1�xu����u�J��>J�翍��0��a�>Y]$�ט��Z�����CI\�[Uh����|ϐ��N��<OJ2�cY�,5K�ʑ�u�4p���c�����H��G��E��S�7B�K3S�*��e��l]	����Bp�;m�V9�4�b�L�L/@���N*��jܡ6Y%Jm�{��ga�gJ�4#�}�t�,G�ql�>�(}n�a\Nr?�93�:�
�,��$ip�ޤ^��=������$z���@ ���H��sv%�,�hU
� ����(�y�7�}
!�ɘD�.NF��$K���h@o4&#�!���Q�B�v��ͨ���58�%*P�(�7�Z���0��nw�W��@"�~���)�zg �j'�@��d�+�k#x���!�(��b��J���S=��0L�t=�4!3���3q<f�%w(���tg��N�1T�5w^��{�i� ��UFw��=������_�c��a����>2m�om���0�H��֠|���k�hü��cg��s1 a�;��v�����\��a\AyfK���
C�e�:��=A���2rAp?ҹW���H]n'm"�yq��=���*����<�~�.+l��ѩ>>H�\�x@̨�
l?�"�ͅY���牬�F��/����O���9XJ`*����c�V�a����L�c�Lڙ_�`h%�g�f?���⡹��K�a�a�:$�Tv�.�Aτc��~b5�7���ѫN�c'	���OH�V���5Xt�Ƀf?�:��_����HM��j���=�%����/�.`�#�X�h�yۧ�p��iC�Uؚ\�G�V����=)�.�[3���/�Y���t��q���9q8!bd]q���P	���7]<q�c['S�c�?pf�r�����ȩ���ڑ�=�z�������T�Ҍ��|���?��Ә���	Ҍ(�K;Ը�[ ^����C?x���$a���s	��M�U��C\�"�t�/e�t�-=��n�h���BU��Jpܢ�Ͱ�����95KgG31��nS}�C�i���!קPԒ�c�cAԄB�u�+JZ x
[���e���oRs�����3��Re�*��aD������фt��:��(������|��.��n��K5��s�z�?^�N[���R�^��_@YP�,c�����j�@��Έ߼�&��*:��c������X��+䵈��L{�R?ӛO�V��7|I�ѣ�O�y���S�:Kc#lȨSK%6���-�vGNZ,ˌ�a�LC����!�fU�/�mo{�%���.q�hY߯V�TV���}
��Kk!C�Ekr����}��k�H�`ⶨ�^�7��X�	Z&H�LT^��o;���,��J46���Pwh�L
��7����KpiT{EJ��;���B|h+�<L��� 9s�AS�1�h��l��;#ء���2�'N�����ߍ�H��lW���)5BLPǣ��IE1������ ��-����9d���H 1Q���Nk0�PҢ��҉��P{��.�]����b�M�q�/=�����^bT�U*U-���7����/(�ŹߋP�� ��ł�! @��}���aW�T�X�gu� �j����ȇ�Zfp��q�/:��n����]�����a|8�d�rG���2�3����9	5�1M���_�&�]�v�z�j��fRtXM0��i�3pa����:�b"��N�@"x��� �+�w�)�>x�t��#���4��Hˍ�kU�1dG�~�����9����[�R��2�6�H3�_tǎ��7���K�*�\o�>1�4���,;)E�(Kߍ���U3�@�����Z�sƥMel�ۧ�ܘ�߱����u����my6�,���A|����Ue�`,��{�8��;��������sCV0mU9�&p�`KF�"�B����s[�Q�:S��ȷ��[��ȧ'���/�-d�������}4\9{�n/��I�_=!SߑmC06�Eo�,���͏W�0Ұ�ʹ�g�|d&(����_Ƀ�,
��9}y6��*LS%6�̓?�j�Վu�T�#Ig�q�׳w��-s���c�R�b��R6�N	�ċ`�6�hg��d�[�~sŸ\	K~ޣU_�Z�{�u ��|/�4���ƷP�f-m�� �\���Y��-Y�;U�5�Čv���4(�-�_5ϾKq��`������5�$iŸ�;�l���S&V�p/�����/���O8��ќ�Blo�Ϭ�`72��6ٿ�*E����w��� �.�Z�������=����(>>ʗ�J�Au��\�B���^fG��G�4{�_�e��: #Ѕg��zp׃(r����pOv�k��xی�zg?��4H��[J�^��~�p-xW��-��Tp\}S$�'��*�=W@�T��S���&�ä%!���@���+�-Hs��祤�o�W�ؽWG��Fv)e�W�����̣����n?�����o$9�R��^CM���YeP�K%�Z��b��[���K���6���
�ݡ����b�	ʓ�ye����q"��A�cǰ�7�FEj����$70� /��_�.(��ҟ���QZ�&d����2�Y9�eob�}'������&��Q9^�
�4��l�-�C���?���;mB3����xS&�~q�ʼ;#a�T�Z��!�� ��-xn������p��U-ҙ�n�d��]�����+�X�.���g��R�*؇CخV��S���7�G}����?v�!��,��_��Cjd�Ӥ����Bb��DGKƞ�̗Gyq���Q�T���ǩ���Q���w�bo+��Si�n����:YI�"�wc�����'�� �S˖�4��V����/ӯ�i�*O)�E�mϋ�K���^��.@�&V�aLH8�H)�L�S��g�j`sb�@���a\_�Ս ��{!��^�g)��Ñ�f#�G���Cu^�~A�w�o!6��vr�r�)c�\����2��9Rm#���=ֈ������_A�DQ��\�����5cm�S-*�����f�&7BV��r��	c�  u.(��tCJ\�5;�� ��ߥ�XB�(cg���к!j�/��4_V���D�!�����}��dԟ���%���^P�L�e���������l\�ҍ�|���:
�F)�+_�r��B�����;cBW�0�%΂>v�Y!0K�kq5���)N���9}�vb̿�M���,a;S�tj^�8�Y�e�����o%�.���AL�g��D3�[�p>BT˹vBd�D{h���a@��>����+6��k�#Q{ �<M)�I���<3X���l�ї�o�[Z��)���]�cA�u�@ò��(')۽w�A���� Ç��1=�{�N���(�>_8�zz���QCT��?�w�#�i��"�������j �Y\q�
:LT#��lWe�|!"��^����J�wJ\WՀ`�)RQ��\~�.���/G�'�����#�)5��ۧ��v�]��p�����]4S���2�4SZ4��Awc���ͷxJ(���^��"�d�����.��
�*�\,�U)�i���>�ɗ�,���T�x��&�v��86���F�4X�?�v��lh�o�%.�׬�m�`Y���R!:{����ǅ��?��v����6�Ʉ�DcX�ʾ�/�L��~ЪXr�U�OW����A�"�K C�s�yrk^Yc�-Z)�ڃh<��zB�G�a%#����z�%�bɅ�3D���.�T�ΜRhmSAt�ߴ�6�'Yl3<tB�Մ��1~g9�e�!�}h<�Hk�'�ʥ����l�Vي��bG�k��9'!|���b���a��?�4Z��E�]��ٱƍ� �r�����LΫ�/\��l��pO�hԡ"H�z^q�K���K���c0����(�/~��?��.!ʕ�!0��U�p��/b�A�ӳ����Ĩ�	��t����q����#!�	D��2�������<p�-X��X�ǭM����x���F��Z��Ӆ���!��u��������c$x�0�1�A��qvQ#D�Sc�'3l�*�h�L���/�@��U��g5�o:PI��HN�0ƪ����h�:F��=OLyX%�N"�S�u����3���{�w�B[M�E� #aq�ІJ?3�ϏY6}��5��@�˔�4�@ji��p2ٲ��ۼ��6ٴ*���ݮܶ�vv.�T�Ng�!�Dw���`?s�.��rf�����My����<�mC�l�T(��u@��5�����ג
C]�D���֝��IښF.(J��j����S��5�u��y�5
�/%*���1�wcR
�[�뒤�%�%'��~��d{�C�y[s����c�O�+I�	G~3�Ch�Q18���Ŏ@�s4����&�+�.#�0%����ex[I�E�g����h&Q+�TDd7�S���$��F�|ȢЯ� ��vzL���q�؉a\���U��_�F#��L=�Pt`z�v��������9rM�X�h���e��"�C�5��� o�,�a�"���]0Ξ�b"5��y�h�Z��E�q����x�cČ��/d�d��mӔb$�q��3ԗx�o�{)�>�����W��p&3����&-Pf�N����LA}qݤ#�[WR�%lh�Fsmͥ�r�2@��t������M�
}84n��6�.7��fl���@��'�^F�|��s���G��A�eҦs`ž�E>t}��{m�@���7À�����X�����G��I�N7��Pt�k�ތ֊�\��[���lď�4~��Z|������ņ_�&/R��� s����Q�މ�~��Nx�_����>��Q���y��Ug:�X3#���Y�?r��������د#l���.O�h�:�޲��ux��Y���>y'b��ދ��u�H�_�<��i�M/C��X-Y�^����OCe�.i]���k�v(���0��uT`o�}Q�;SˌPT]��e��o<B�D���;�y\[�Z��F� ��?}�ô�&U��� �L݆%�9�H��G4^���L�%�z���� ����'���H�@��la�S[?��J�@ɞ.�}���A5)=�P񋪖0�(_=(�N��S�qŁ*t�P�Jy���]^�CՒ�%^�[Z�0�mA^2��{D�<�U�X�Ӣ�G�s,z	�ߊ���`(�����}�z�P�����Q��l&q�����H�~�1��cf,���pCfá�چXN�)�B���u�2�l�+Q;�����'�a�^OK0��Yz-T�0�r�	pCO���B�Z���z7>��7i��'=����2�߅^7|�3�O���ܺC ��OWYDe�8�ތ�x�DQ V�Q~-! ���EC%W����2�O�Z�i��tq���U���qv��L�7� 6/Ug�$�9rh��*ZA~R\�'�[���#w�*�X��<l6�L�Xy���̠lc�Lv1�Z�j�C�2;�Aq�	����̹���9_����IZ^#�*
oQ����ʺ�:�L��dT��
[�j_�S�scT����T�h)G\ewJ+^@Oe����6&	<��/��$I#-i���D
�+� Y O�'9CnoD�V�Y[	�e	�}�����p���a�ߠ����z����~@J'[À�;�!�#���Y�Po�Ef?�e~�ܰ�p�TDLh\�oЧ-PO��t8t����Ãht���	z�)�]�S6�}k ��+T��U4:]�Dw�lÄ��jǏ��NC��=�\B| <����s%��,~���d�9̒������;��Z ��0bj�f��
QZ6�+�ӼhJ�Nvfڨ�H	�¨T�r��T���T����EH_7y�G��|�C}K�d���::.ߴ{I�鯯�:�&�u�[T���L��_/��;�Ns
�h�h���\yQ�_evN�C�
%���A����߼��뷈)��lK��	��6<
X���2 ���:��f�N���K����fӂS�|LB��n�k��@_ד:=V�q$����;Vc7�z�y����Nm�`;o�S�'.��n:+���Y21�H�W�|��A�(�K��-��*�3`�%�
�\J�D-U�LR4Sc-��G0��y@+>`Ba�d�y29l/;$����oh��~�����*
��L�񏷍c��m��X��>�d۷B�zr��:��@_���g��Bʇh'�C���8n�"o�U�-c�[�u돬��DM�l}�	����o�3B^�<��p\�zE�t׻�y�{bq®��ڽt�^�����,Ƀq�'�Y�<ɾ���Ǖ���V��3�&��\�(��p+X�<��s\A�!oEN�́9p1��0vǿ��8O����㐏�\8���;}��0>>����ꌠ *rU"xt�j���AZ��oc��~,��8�|�J�hub��n�/���� ��ŶOCg~%���K�{N?�o}�gNfI����M�V�� H���)�w��c��U-�ڸb��N<Z����+2LG��t0�i�^š��L����S��<P�:5e�zm�o_�,$*��B%/��
����͎{^sqLi@��
�G��ԕEߥ��L�����.8��G��
[��-ݾ�I�cŻ}���<:�h���ھ��S���q���u�����4����ۊaV���������
��7(�)X��O�St��g���qA�Н�T�[��4M$t��<��
�b�ޚ)v�y��IR|{��k���m�1�W#� ����͐����,�h��R��SN�����c����yA!�#!r:����l�+�����B@nƅT6�YAZ%+j��v�����l-V�����~��� ��1�mƧ�Ԃu��V���O9P�,6�v����Y��"�q'(�Nn���(��Ȉ�.����跩��_��S��	ځ�;�H�
ţ��8��� y��1j�$���������"R<�@��2���Q������_k��%������=�ޫ�;�)@��ei�5��z*;"O�M�?�\2;�m�/0M2MPDվ�H�������gk-��m��֪=��(K�6�n�4��՜Eٍ��X�2������x��_A�1��sq��R$���SO������(�����#r��I��A%�������>�ȊH#b�P�yEH��~��F�ˀl&���1�+�1b˸cB{SϾ��ٛs�������ፙ�Y�%���:����`G����b@���lЖ�7����0�l�D��;ʳ�`Z�aX�R6����6�9K�����6���Ry��;ۭ/g�ߕ�����0�.�7)�K�~�������t�����e�P�O�?��o�4��O���u�
��^Х; @���դ23ޠ&Z��� �7m�m�q*���\��&�-�~�=쉏�ק���y?�˷o[aS��)׌�jeG~�,專/��N)�y�����b'E���<��W>���q<�3ىm�������D�����(]�-g߭Aƺ��w�A�!s:����7''�
hj甊��5;�3�3%��0L����wYQ��x��Oe�{��3���_���ug�g	�eJ��[��^�rV��/o����1�!ǦD2�:����Uy�3A�O�PhV�����?(�/PG�ہ�KZ&���~<#��˘>
(�`K g@�V�_Zb�q�ǋ�R-���`�����\{�S^��Up���c
4�B;B�[��ym.�U���x~�N0K���\V�g3U!�?ߋb��n!rn0��-���6���`�L�y�%T^Z�9�q�}V�5软�~���+�*�r[J�9�m�������@}B'>J�Z
�B_�i� e�NP�l��8H�Qh:[��_��������A�!�4�l���2���4"��ES��y��ع.��Q���)��L����T���%TS�Җ���Ї_�\Wv�����'�O�Ǆ=�'ޕ���jh��u��̒�9g\F�y�LC�ʝ/��Ax-�	W���`��t3�i���d���ASD���e]�"�y/,r�9��]����D�� �MH���+�WI�>V��R��Lu�2;�m̥�(�P��� u�D�������B�Rcٙ~�e�A[]���4?�vuLb�UZ�P��1�2y�Fx��حɮ���@%&/C���9#�3_'��[ø3�<����#�����B٪�G����u�I�W�<�@�+A�����;���Ɂ� ����Vj�����?!�d�n��Jka����Z,�NTkaU��M����sbf3&���nmNE����!��4��{a����꘻J��Pl��7�Y�ӧ�Yd'_�H�jph�?q=��OZ�f��[A+�H�Y��u5��̂����u�c梣kv�F�>H��D/����9ڌ\�E�1Ŗdh��V����k�d���n1�W%|I-�����H�B�������C��jʈm(��IXE���Ԓ�D>��5<6�a㝀����O��r)�Jk����B�g\u���2cs���@��VD�ڒT�A
�P�s��~�;�>���w�$-~���ɗ��6#L��$�R���%d5`��iy�o&�}[�/��c�o�8�kk�r��|<�Ҏ&)ݏ\$�Xb�a������J}k$3�2z���0e,��ѧ(7��㨭V85���Ez<�Z���yߺ�=#q�"�N�2��f
 �/���=@��L�)a4��ʀ,��G���RX
h��~-S�7.��b���J���8Z5��ب��{�#�	 ��d�2j�

괬�z娱ρ��{�˱^Yx3�[�U�K�eR[�ǤU��p� �S;��7��"�h��/�_�6��y�st��Zk�-��>�.',�Z�3��gs r��]_N9g��4�z�Uu��^L����!�U^���iEH@�#`*i�*w�1���3�G`��b�E~p�o|�G�����lաN�<|A�3dPiig��5?��Q��m>,�}`F�(��Oۺ�����f�f.�|�I`;J7Ac	z�񙗷~&q.JI9��cj��W�A�p�0m����/�ޯ���.A�͞
,�7����
}�C��q�oO�3ȩH�f�L~�����z%8�������Nm)���= ��z<��,��?:$6�K�%x��;m[I���EZ��;�'S��j��vQ�n����Z� �B#��ű\����~«��E:j��Ae�ң�
�d��`m�ԑ�n����<�)�5�V$�/0�o5���/�Y&��^1WR�'Q�UY+>]C-M��ٰ(o��:���KЩk��	����~�v�Uja�5���M����I�	�mV⧦�MXG%�"��F�� Y���]�n_�w�r,{V�u��NQOH���6�}�WNt�c"m��eL������G8�<ME7����ƥ[�2SHQxL��C�`뗁�޶��RB*�7u�pd,�
�"zTp�J�NK�����[H'񢝾P�XZ�zt��1l�%! w�2��%.�r���-7�$�4�s 7�iu��7K;���`%g�����D�	�q@��|��3t���ב�yZ1"���yl��W*��H1u)��](���V���R��5a�g��O �����#�5s
�ϫ��<����S�ٸ��@�
B�w{}ͥdmh����ؓ�;b�H�)]%1�7�rI�~��`ə���EסA� j�p�N�W��L"d��;�צ�?��:`\V~�z�7!`	j�l�M�3Q��ЖW!�vBʻP�=��,?&�P��|�ro��)5�yU9�l&�7��,�A���t�	@�}r��'�(
l9룔��n�e�C� K/i9����� L�v�&����\�ʉ��>/(�?ݏ��m�	�y����L;��o0e�/���)�~���_���Z���4�EЕ��B<��w��Hi �u57׍mO)8��Kh���n��~�2���;������G��~���W��@a� *H�t':�xC[�f�� �.����� ���w��|�{u�t=�:l�px�Pq��t�w�j<�|��@�eH��X�Q���+�2_W��Ŭ���KR���#x�x��ԇ�l��h�4�ŭ���F)�����roqag0��X:���v���j�"�~�v�5�.B�g^��̨9�!�Ч�����DS$�R��m�qU�orb�_P�]�ǌɏ�
?��ԑH��yO����5�l�:����)��T����/P1`3��y��B(n����*Uxmlr��Q�+v{7d����_da�k��`g��D�O�I*7%;��-;�ۦ�2��i����o��.ӑ����a�hek=������i�9]��[�xT��3�mmL�3s�Y�<�������?28Hc�8���<��C9V�@ſ�ɃE����>l��O��[�00�Ǚ�?|���Db���P5�s:�E�*E����i�2�!�4!��p�Ł�}�y�0�F��hd�oI��@�X�CV��*�p�_3e٤��;�P�a�jB�.��&��U����f�tIgL��"޳f꩜R����ZB�����C�V��U��i�K|u�� ����Ϥ��V}GÞ���Τ��!���tK5:[�α��H�`y�IL���ak9as�`�U��Ƃ��.����$�J:2�&�7)W�GrX/��S_�'� Cq�#��T1Eg<�)˝	�v&#�����������#=.9ٯ�;z"���E����e�MhM�����KOL1(�vx3����������������צT��z�Q��Zaǖ��HshRhn~`Q��J��EM�2}�lɏ��+���
�%R�b� �$V� �U���k
�}'RZ�ά��l���$&:>=���~(����|��K=E�*$;�1�`�3�!'h�H:���ƚoRӜOM#���q.$���"���� ^Wb��#�&�0
�x�"�����pd�ř�Ba �/rIB��.q�^���vG|D3����~�Վ`�m��afb�!�W=@�'Gz��n�Q����N�R��Z���@��dͲV/�@%��n;��{0�����a4!�!�H+`�F��v��`�⟬�24�f':p;U���a�s ϖ�s�4���+�'��(��J�"	%�W�9���d.��g���aG����OV�k�'����1jwigD���N�M�y�=n�������^"h��g3����,i�nP.���%����v��V�"z��CH��VXtAqP�#�qnv�	+GG.��_ ��bX5�bN麂�����BD9Ktj9������Z��@y~;-��IQ�:J�ĭd9�N��yk���{�X}A���^��'��g�ҙ�JT� G���դ�ڿ�����A
�`!	�u$ؙ�E=�P�MZ���"ŹK f7t%�|��˥�q"@Q��b�HOK��j�!��S�����P�*{�B��:(\��Q��I�І��s��]A�����B���Ճ�},M�M�Ԥ��5F{8�G"���^�������gL�#W���������s4�z�I'����p��OM���|�g0ف�%e�c�_�E�C�]���|�;�Mv�M�@�_��'�SF�(I�d�({�6�����w
�|E\g�"�0F��/�7"�k�u�$mvJk��R�-.v��G�;�֋|< ����)4f��M��y��7rv�3��G16q��E�5���G��R�nB�sH����z�@���z��O�|�<��3�R��%� w��a�ۑ�Q��mb�op��&#hI�P�'1���a�5׼;��2᭘�jtYW�7�`[�_����oX��9\P\1B�Θ��q&�h[]�� -ݚ0��0m߼$��<s֫be����'���e��ǟ4{�x|�Q�^0I_x!��譓3U����~G���W��ɓ���j@&zJ�Ѭj�ʊgW����K�3����s3�;���С�n3B?x�焏L����?6�K�(�1�ۯ����U���DZQ�%�3+��Q�FKs/B�n{�<S@V!*d��,�z��3/F8��<:��F����7�X>�n5���sF
hSC9z�R"�$9U����͊C9���QtL0{O.��*�"8"	�n pɞa�〕%��2_���4��M�5�n�F����%���� ��1�5 �=7��f�LD������}��8=��M�^�$��.a�|���CYA�o��0�.L��f�q_h��M���������L��Q��z.��QHJ�4�[?��+C�'W�`�Z:r���0�YP�]�zN8�x��p�x��)�h+���,��;g�_�T>4.6G��
�����u,�ZK�����X�([x#�?�*(�c]OC�:�8������x���F�>��Z�a�V���"��m��^_��q
�����&�↯s�+�g��]kI��s�ۓ�ڹ�&b��-赟��/'��xr���i��?��"%�<ϱR��Wr��3c�=��Ju���ʕTɒ*��X6���E�W9��z�Z�H�bt��0�:�9+J*�O��$�H��Q���[D3	���"�A�?�4��Q��s��J�~��\�e\YЬ7�Ν.�+�Lb�E�]�(tCe��5a�!?ޡ�PrJ�f�bP]����r�"ƺ{g�a����r�;���v�ZB�7̧�Ad����H:��50[T�?�덠�_p昮�1O*(>De�g��%s�Ѽ^E��>\"	�⭋�-鬘������L����(b`^Ew�KK�u���AIS�}�Zf��G���/�*ՙ��A��.�F[����av��E�=��7�r�Uu���ܽlH�ٗ��;
�iV;ѹ��5�R�v5��b�+�p���ig9���}���`���%�x��s�q;VJ/�=��v�4L'����f���yH��a��VW�9s���~�.��Ғ�/����ό��q�����?4<�����Yܗ�Sx�1��N�X�����3�������`J��������!i��[ȿŽ�]�q֦� �9�b��8��A��{�'_����4�j	�:ۋ�~?�awZZ����
Y櫉�A���DW���0'ҋ��vB>�yMī���O�)�鎷t�(��&?���%�L�	"�X�`*�D��a~�N׳�O�v��LB�,��К�uI��� �����<��ƌ~x�@�A���k9�am0(B�7K��j��5����8�k������;�	�����;W��Y�p������~)���c�
oCf����䑍Y��'ةTvf6���i��@!��cw����3�(�� m�GE����^4jkڻe�x@�-�}�ބ�<&�L֓p$�V�p�A��f���4������)��9�tW�a�Q��ݩ�����<à��Kq���.�ԕ51�4튦����G )�	���j��%/���҇���-�züO�ѵfz.�
�l �bi9��>@�D���w9�d���6��f�+��/iH�^���ܸ���-ړ��X/�x�L��]��1l+�L��E��u5�(�42.�{��
0 ybgz�1��"����m�a���$���<>�O�D�q(����F��qm�yF]v��|(<F��$�]���.��S-��ݏ���������"�-��$��q4oH�<ػѦ�Sƪ��+���4Ź���{���
5@��v\��㌺����[�[�st��e!�I#�}�-eGC��gl�ljbZ���$��S�6P�%U�ZL�M��E_C��I`��;��خ9�%#�x�~�&�=��r���J�h�~�S�Ѕ����?<A�n�5n=��щ�G��c��5)��BQ���֎�\��b�ۻ1Ggj�>��bw�E��I�UVޓ/V�O��(�����fw�x��Sx�t�Yx��n8���?�9�+(����z
���1(P����ɩ��#��)��tPc"ƻ:�4j.��(���+G�"yݺ�ek��EȳVɓ��Rq]�[��������[Xv������I��.��y{��#����$�_u	Hu��g~��K��V����߄x������W��`�i�k���+ф�K���	�wI?�rs(t[�(��[���Q�j�]��9����?������C[(�!&���[�&��[��#��R������h�����t4k��!nc�
ce�ɓAԣTa����T��Ar�~b8�V#~�7�)!6�m,�$q8��U�L�ȋ�Ǆt��Sf@�/�E/���'�)�{S&�N�/줳�m
Q�����4���u�O�}b��S���m�
ּ�7��=�x�7i6kf��"N�,�54�/�]��c9�φE�Â�]��2J?#`a^\ۙW���D�T�x:��0��C�Ҵfc�D.�Ui�A���C�p�O�ɛ?�;Ô4����ܓ��5��� ��ߥ\�� )7� @%������Y��O-bw�( �'{5�����Iw���q�@t%ɳA�~1�1j;�
H g�ӳ��ۨ�y�aˉ���矆̕�M�Yl=2�Z��R�-��ʎ��Q�="�f��%P�l� rj��MJ���lZ�S���eG�J&����!V`��k�M���SH�ؿ�J?:Uc������=���C�Nxb���[���i�����ԾhL���K�{��p6�������(��v7�v#��y��j����&���y�0��˩m���z�ٳ�9���{Jd��Ov塻z:;����'��6pb�NN�5�g��`'�*��T��gBcĦk�W.��)�x�����q�K��+�;'���Q�U!��fW%J�=����=���|"&��	����F��������������d��#'�޿�K���.�h˷��,z����'CI�x���S���zi��h/n��:1�;Ԩ+pz��)þL��ݙ��m��T!S�K<ڍ���>�<Tx.��TFȄ̒�WBj�f;�>��_G�Vk��-e�P)`B6VF�X����J�L>ob}Pb">ы�$�ԉ�
��Ը�F��m����"��Ӂ��mߧ���%�!�P���-������V�Sc��p�*æ���ߥPc�XS�Ȧ}P�㈵��o-[2���H
�uپ��;>4�-x��i5�7eg��A;�v��X���LK������q��ϒ�8�Lw��d���Ul��D>�O��!����Fɟ թ�D�̸�z����Es�gU�ז, ���6n!/=�U�h�m.�s|<!B���Q,��>��$��^��@�g�j���h=�/���s�~k�kI�LKwq�m�e��G�w�o�l�}�R�w��_f��L��7é�8����s{�99. C6a���>��qԌ"k�@~����s��3�z�4T�K��q�/�8�Ζ���	���**m�<rϑ�K��f+��  ��/`C.k����%/ߚJOG1|��
����M����/�����Or�i�J�\͍D@3���?��ʖ�+i���u�A������ĺ�c�@�?_s�o��	x6a�7H��&, ��v*�ۗ0L���j'��q_C�2�],�5;���$.I����.pܧ�F~�M<��[#$ҥu��Gr����J�hȽ�R���PV���&��א�_q�x<�sޝb��� �����?��u�qo�Q)�c�����t�`��0�n��2M}p��mꈒ�ld����S���X�&G����F��$9̾+oǠQF���A��귳1�4�?���x4t~U^߸\'�|����$.%�+�� �'>q�t\���1��O���Q.nn{ĉt���A�YΞl�m՚B�������D��2?��5�b`ԣ���世(E�yW�hq�]v����~��9ы?}9,q�w#�?����x�}�!�5ׯэ����A�!��$�|gN��y��%�O��6�XHT�n�0��?T}U�C0�;҄ذ\,s��Y4��}��#Q0A���������+��N��@�:򺤃��譆��!��\
��l���`�q�d�wJV˯�JsJ=v|�N�3-�N��(~�	�/���.Gd���s��&yn�� x����)'�	A��@�d��z9�H���vy��]��څP܈:���$]�J,�ؼJ���G���7�� ���&� Z�C��4SāPH���te}�ĀF�4IןC|L���c.p�!�O�ZH���ƙ`?QS.L�v%����/��O{In�QnU	Eϛ��0v[����n�/+�m9�-�Ӟ\��y��(:|5S��_/�X��dK��?���ư,3�nڨ�4����j$T�we�Bn{M.�<�T2T�I�Vx��~�,W�T �<�/�)���3C����Ǳ@$u���[8
��u����߬q�ˀ������ �Ƃ�h�p�:RkIFY1JY �+�Dr�P:���&"k�@����;����wM�sST�!R3p�{�o_���u��X�]8�W㥢rQ�V�ih�2�H�d�8�
ӌ`BE2��G%>l���}%�b�ե�
�q���)����r�pZJ��e���Ļ�%�lkw�Y�ɼMY��4�r����P����]�-��F��3a��S\Ä�<�O߶���´be��9w�k�
�o�Gʭ �5���x�
�KmoD슭���HV�� ���5Βr
S
6����; ȋ>{c����&طڲ�~��5э�5�����.bv�e$�٨�krF�Rn��R����T�B�/%�!��~n$6��w�>K�J|!�R�3�ɜ���yj����w����G�����N]���5ץ�B�q���˲%��H��Y\�|���юn��%�(=&�����q�2��)��q�C
y�/���x�����1�-7#CO$�d�����Y[���d#�|��E���og2N/Oޭڿ݇��ʦX����-Z�wW�dI3��2�}N,c� Up�x!"� 4��!C��
�!y��ڱ6�3�?�����II�j�Oz,X�"��6E}H��R�Ӫvv��xt���A������Ӎ>z�.:6�R<F�J��&��0Cuc�����ճ"r��z�q�0R�:��B�N���SpCR'���Z���k�`��`%0���{^�*�iO��5�����jܸ�̂�g-��}�]����N�5��&l�?b���� ߼����Hyx��M�Q�&{�X�l����S�������8#Y"�J�3�;���h�����ycK�5i!
�)�R|��圵��������,iKc�}��$ͳ�cؗ{�_��@}����e֏b��1�=q�5mxC�F�/�2����c�ᙷ��:���B�4�g�?��1QvF�)��G�B|O�_ y�'�X[ԣP�f��b�S�����hF���g�uôM'o���Y��m�9��tsX�I�����qkyϭ�bn@Te8:`�>��m�p!����l����n̊��rƷ�O�8C�@��w�~T�҄�1s� �$�減����:[�=���ُ�ܜ��g��Q���_O����
�Hy���*%M|v��cm.\�w)еM HR&��T�xZ��D��"
�KZ)l�9��.8�cW�3�Eaxt��d�n%'�8���U�W��t$�6�8 oG�b��ˠa���V��c�1 ��@�Ӻ�D�}|�`���$�a��(�4�y����3p���G�L�/.��V��P�]���o�+]	���ɱ�qnb@$>�^)��Ԝ95ܞ��o�ir������G�7FA� ��k�L������r�)�"��ȿ�ZX�,��]J`���{[ٶ�xkSk�����͹��:����JL�]�=s�������ʸ��l��ߥ%���b��_�;�ك��M<�|ɹL�eO�����\������4�c�P�U_��vw���:26�}�E�5U$J���XU67��+?sZU�`�ݺ�*V�q��$L�%L�kL"ÙuHf���UA,e4���	�Q~��En�0(:"�� ��S�갮1>E�i�g�T[�7	�Lz�����:����A�l��P�`~�o��o6͗]z���m���wR� [j��g!OȖ��KK5G����˻8�n�؛͋�OE��CXƺ���O�V޾1�FѸ�TI��ç��yt�/r��Wq_A%xId^F"y�������Hx����yT�/V������vPlu�cߞE�V��Jr�@<=�>���QO�sc�:K1K��^~�	PZ-�z��>� 7�HK1C�׭(�-���|�7�B؎��=��p�x��1�b�1ʱ`	�x2���4$�Y��{�q$g`ן'��E~O|>�C� v�b�o��~�Xa<�.�	�^����O�t�I�!44p��7�>�R5,_���5�5��A���e�S~B�,r����hb/�6u�x��ļ94ˁ'2�(5L�O�g�?���NI�'�x��U�3э������i3��1X%�����M�7��ӄI�Y[�:�	>���0���«`a|BbϞN��Lݸ���{���&o�5#a�{��z����'$:|iU�pZ���X�ݤp�62�k��k��;��-njtb �g9�)7�k%�~��9qvz.FC%@_hvH����#��d�eN9���
��x@�~XoL�?��;.��	8�����G6�������y�v�0v(34|G}[�njAKt��2_/�2t��X&a�a	4�FB�W|P7�Sh1��4���.�E`�*����fOۺ�][w�e������ۘ���P1;����+d��״.&{T��)�q~�=Z��n{�7#dDϙMEC肬��B�و���+E�e���y���ul)J�%v�9��{�=�>��'����<�B���-K`#���02k)�V�WYR
;v�"z0���x'�;��dk��'C�m�e�Ћ:U��zh��R�"sX�fB�6L
�6`��Fm:">7��3���7�(�w�#�q��]��$��s�5�(s_c���⿳�\�<���G�i[�Ŀ��tY�����!l*k�^��`y��ߡ��6���/����~H<?��]�8�8d;�t�$�5�&�]��,�5K|K�����ߎZC}��@�kP������f��Ҥ�><�����_��#��v��
��A��g�p�rTx�����-�;��e�	�+��������$�/@����"a����x!�;�UvP<a��&Ar��ɬ"�^��/wkkV���=*Ԁҩ�-?�Ͽ�/�*J\�J3Qգ/�>؝/0FŖ����U���68=v_)*Jr��]m�Ut�����l`����*�v:>���&f��P�aV�dKq��?�`� ?���u��m[������>q�?,��������u��vY�H�aي2��}��~ `�<��<�ۄ4˂��hL%����k-��AS"{+��;:CB�s��Ȫ�P=�������l��z�΀v�! �\�ʎ�W�<�}.�uGZ����Z.��h�3��v���>O�4��Rّ�����i�Z�^I�>�$�������*	U�K�=a�$,w��74\Xݷfx�wN?�K����8<���M��gb�D�t�<EL%w"�`.Q���nꦈ�G�=��]�XB�a�L�_e?؛������EZtD���P&����������K�:}�
��!���V�#ΰ����3��@�T�9��g�-�(D�;ۨVP��lo����=��M�^�ٿ��dqCc<����Dm��`�y;�Y;1҄�r8.T�l�M������̊���8.7Izd���i��Ě���9�ح��IT�G{"HwH^*���`	�󵄍%W$�?\��{w�l��谴_j|"�?�O�A9jZ�Iq���C0s��X��cM�O<��|� �@@�3�͒�|�B��j�"k�x޻N"��ʍj�ǵ�E�� /��-�*{�Q�����|�w�@�ӗ�m�$v3
��xw>��y�C��n7S�k�l}�8�p?.~�����3M��׵��ců
���N��N� 	�!$I���M[UL��~l}$CU��ĩ���E�N���-��Cݘ¢��:����{�pB����4�6=�t�qS,W�B����a���&'<��5a��ׄ8������Nh����X;7|��:��Bf��.~��o�z��?�d��]��=�hN(�T3[ uHF�O�[����Tp0���*@ x���"�n�VK�,ȭ#MI�%1��0�1�j��� 
���3cyZ*�|���R*srO|7�zXB@�&�tJ�H��+����/IrC:�~�Dej�f�"g�E�6�0݅��XuC�c���>�0/�)+l���v��U��Ad��[(�f�H���)gm���U�-i&c_l���J��b��m��T�{�.��ʑ9P�4!�����.�]/-exIp�erg�^��w=�$H�D��<�dvl��ӤLwJ%��eT��pK��Qn�fq4m���vAC\B -�����}6�#�aWQ��54��x=mVu�&���"���vw�^8���eMU� �R�����6��m�ͼ]�(O�|�0M�&�����f���G�,`;�ez%�WF|j�%Yޯ5��b������xi�;㧠(!�3�
p�U�T��]d}�0�;�����QÃ�X�[��JC{��p�ܬ�uҴ7P�q'�,�����k��'4��ҵE��Y����$��҅x�W�'\b�>U��֖<��=��#wSԎ�7���o��`�\�ي�L�^{�E'kJ,$�[K�=[�8�D��wwB��ʄ��ʵ%�@����+{/3	��{�1�oӶ��7'$dXwL���uf �u���u&wR-Dk�27��¦6�]�F!ѱdx���e�=Qo��i[�2�x����D�x���3թ�_�f˒{Z&���$����h=�Y�B�5j,�ӌ�#WL����0H1�S�%P�!6�9qh��/R�ʒ[���Jn�2�����G���*Zb�Qj�jM^m3�����us���h�Nk�!%�U/���YA&P�����O���gC�6q=7��U�D8cYK8u}Ў��7]]��2+�f��
,�h�'3���ʆ���BTx,���6Y��6U�yg�	��&�
"��L�HvC�X<aS���1��]F�C��<�WeL#y�F	�uwd'�2��~bq��z�]�\�p����VY�f@P�3��kNy����Y���`'
2��w�on̩t�7��TX��7n�`�m���8���f�x�˼�k���?3@��	�} ��J�g/+H��}���/��n��0s�%�V�b��{Hy�T��m��=0��=s���eEiҸ~ǳ7�@�$.�m7�����2RKEH���<������A�쎤҇fH�v�F�E���tK�H}��Ra݅����?�U�-��ڜ�� ~�=�h��/d��{�:�ɖ��ړ��Zz�9�Q��Ub����9�8�Df�bu�3���J�u3N܀z�� �
�7L8����������������R<��԰ri +�T�k�y�܍����hjtc�5Ffe����e��|�PH-����b�C7d��qAB����D*�J��o�c����1|ͥ����	3�Y,*p	9�\����ZXaB������p);r�	ɟ�#i;an��@k�r��{0��=�8��$��a[�U�{g�݅��V��`�m����9�EN$���(�33⢎��}+�oy0������Rad�u�~l�5p��,�b>��R��F���K{�4<b�������f�.���c���V;��x�;�6��Q+Jgf�!>�Gk�2$�:p��X�d��H@��Wh��z���ꦹ��.a����X��<�P������ �7H��5��qU��G�qٟ�jVD�s���/Y���V�ڸ�Xd�vq�:�����̮SG��2""������=��w�"�����5�1+�arÞ&.���(�.2��sq��VɅ#�� e�QKc�G�v�pӷ�Q��(���H�$Ƞ��y��gB�|ݐG����g���k��2�����d��xL�������+���_�R���~�ZB�QT��s�*-���@�)~I.��h����`0}�uTl֎>��X������B<��U�Ttl������Eb�2i�~��PJB�*0:j�i�s�F'��=Q���Z�`���Whq������So�.dn`�#ݽ/�a�@�5Qm%�f�	a��L�"�m�NtEW\JM*�~h7���(���Mۑ�	F�]@��[��&�iy@�t#-��f�������ɧ 3�!ɋ/ݔϒ(�� t��S���؛���@�>����u�����e�R�Ay�f�fߝ}I�R8i��qq��qF�m j���uM�<h;��Ԥ�iXxQ]}�nM#`n�8�5�lf����6�R�Oߣ	�{�d��;�C�&���(��a�A�����pb���7�M^PM椂j��o���C�E�"�˔�bN��aҾ<l�4?���'��:1%�C�)�CJ 8�$O��뽚d���^��C���ڡȔ?�wf"��_�	!Y`)��t�h$�����P���^���3�nhɁї}~�tj���<q0@"�c�j�H��9y�=(��e{/:ܗ��}�k�Uj0➜��C~���
�Ν�S'��VA��+ݖ�)#�%��� �]����r7�xL�F*����.#RKt|��Eqz���U�,�f�}P>�DD�Gj��Pn�2(
�S��J�?�W��"���WX����;�������0!�n`	�������]!��|����������LM��V��y,��<��*���R�@��X鉲i��<�8z���4��[�|�n4j��i����b�`���M�e
������ҧJ��C�����ߍf�Ĉ��")���d��%���dɉ�p��'@J�&�>�b�9裩�OR�FyY��*+:��ɀuoTioȞ�b�Oz�#1��a+�:K5�ߙ@g�/�d��e9�R���R���n�Y������dUY�Rd�$z�oՌ��ϻ�{��[,5���_|�*M.�����"�x��z�����K�J}11�-��H,2E�b�O���á�a��lj������݉`l�$�U�s�a�Q$/=�za��8�P��g[��~��ީ�/!J��j:�K���!ht�4ݎ��9��8�G���:�&T�w��#��+d-;6��nώ���<��r�
����O��١�#l��s���MXu�a�R�ʀT��ܭ����������F�}T�vߦf� Oӯ���i�e��J��
N��滩�Yo�M�Ŷ��L5'�qox<��5��E�Z�&�D87(`9#�_<��|d&�.(?B���W��Ee	6	F�4�_�ro�p<�ƕWm �%=8 ̬�������s 1/����9 GBe��FuB�������~�Z�D�U��u涴��&���m�� �Z�y(�I��'ZB�L�>9m�t[��/XY���w����� ��[��sf�a��� mt ގ���'c]��Q�p��^��=��|{�wM�z{N�Gq���&Χ�U��Ʊ�v �F�@�u�-��r�1NJk��s�;���_n�w��I< �E�t0*G)��'P QͿ�\+�=��돛7��}Թz���J�����l �P`��#���c@��)�Yz�?��;>�
�ϋ�R�>������2���K���;�h؉	TÉ4�Č�&x�ճT���cD%�v"T��9�XA�ٴ5�8#gX�$�}�������&0H�����Eg<�kz)VF�ė����i���6@@�a�Q<�v��:�w	�s��� ��Δ�2���ݧ��� �2:�bzsa�^�''d#s��K��D�!ͥ�V"r0sn{�h���)ti��j֯u`�h�BHΘ�
�����nn��Z��v	�Q�a^��Cy���b\��;]^����9��A��K@W��#s-�U'�k0�u�Izݥ�t�Ħ�&��4N~���&X7�:�{
�3jj���.�9�ݭ��F�!x+m
�� Fv�nh6<��&��!k�Jm3��I�������w�O+�$0�� W�A*��d_
W��;��)�p/�n�t�$����K[�^I؏]�Zޘ�^��Ʉ���@h���h�p�0����^����� |ʛ������tuy���>w2~l��K�
�*8�]dD����Ś�O�(����y�ԑ%�\�;2���t-�6
�m��}j�I~6ܧ�k��g�y��_�������=�>µ�?Zf�nV�!2��On��g0��$�]ԧ�m~��j6汅�߉�d3�<j��#�b{��\�m���wV�ؔQ�&u��T�6>�{�x��-�Q|4��*gē@!9�R�-��t_��UᏂC�s����A�:��0�Bڸ��*$U�u�\���[}��M&����:�6�L�Ni2��T0�|�Zb��Bm+���� ���MiQ�j�)q�p@ƾZb�T(\ �NZ��B��+��P�Hc,56I=a�o��V����D2'=ֶ�b�
专�I`$8k����{Pທ���ښ�ǲ�w3*�>�yMi���\N�F`���VD�!�K���ٚ�Nf�o���j�fB�{06۳�)J����G�ā�Fi��~b���k��\�4,�Ĵ"!�6�ds�s��c�SN��#>s�AeXdl% K<�`֎V��1�7wwM41d_KQ!:-���U��-iO�!6�I	iv���#~���
�T�3
P^~�ʧm��s�_�ϫ3l���,5��7��^�6������8��r8 ����=*O�6��d6�k?�Qu�M̏@��lʺU~��#����弋8�b��6a@���s�wGlI���8�YC��"5!�u��y�qkz��j�蓶�n��

�%G�C�g���(����Ԍ�ӭ��-)�l�cΘk98���@��Υ�%8�L�{���Ï�M�j�@�'�~��R��(BڽXT�y��Y�C �T@;H�Κ6$3s�N�	�+��Z'�*�L=��H��o�E��i�h�M�E�<F�+cl.׊���Z�wp����D�����"��c�����8X�E*�h�^�A�hV�+-zV3m�˻��1DA�\�oċ~����.�H7wv��=&�=����,��EƚBtP�UC#�ɞ8D�(�bS�@0�̮�|�h��h�܃�!�Q[���t���k�5�7�f�A�r��t)�.�� ��T���c�������6>i�$� ��|Z�g8�r��L��YPz�e<���ޗ�b*x��U��E��:��{ y��h��'�&�Z.\. ��V���`�x��J���0��p/�c:k���vw�?���L������'8GZآ�/UHv��`�#7��R��n�O�V^R+�W��'�h[>E~�9,�V_� '��%�l��V)S�Өp��QY��p��H�x�=��$pU���S���/֜��.��<��r��.S���v���A�	�IO�T�y�N�J��:-���q?V/�J�/"ONpljc*Bq]F�� ������z9�ڽ�
0��X��W��b����_i�� �&�u��z��V�g��5����^�p��,|�/�i�9��F��Uȅ0	ۢBp�T�z�;~�ٱ!a�^r�ې4BnDK�G��'{�ڈ����bP�/���B��T?䃰���晡4�,[qK�]Z��[���QɢB2�d�ۜ�mi�u�Rv��2v-�r����C�}���-.��l�5��Ɂ{z~���\+�+�i�zgǎ.�P�2���b����a�õ��D�(�=����ee^���D4��h4y+O�f
�EC�!4&wYӈ�+�cA���������M�l_�ř��$�f���4���>2ܳ�
B��#
9;��y��(z*^���WAuR���b�߿T!�7D��ʦ��������>Kb{�g;��2h'!�#ڪ|T]��Ĝ���7��"[3^��1�L�E��958Sla�;��ڶH��HS��xBd�U��\�É�v_^�{�:zgg\�ǖOrFF�-�%�s��. GѰ�"�hsϟ*ږg�b؛���#;��ܧ����Wo8�����>)9�8�<��-j�?zk�@N�z���������2|�~����+`�#����Hp���I�����']l���b�_n����T���-OΎ���;��� �g��hZ�� La��|
ĸ��Q�GP@^I���س}����5��r�l�m�=���R%�λ��|�z������Ĝ/�;7�V���ٵ.ڶ �v����Qރ�h�;S;�	���ρ�f(e�y����f��6&����RʈeŴ�H=ϚcN��ܮ��p�]��+��A��`�����(�gy1�V����F%�zHik&�ԳZw$RL��d��^�W�RH�D��S#��N���@<��>���]���?��u�|3�]7���)�a(�;��Zͥ^@�.�B�xh�
����8��Ǿ��5[���b�h5�HU��d��3|�FYO�1*�J��f���{qҨ���Ǩ�${S1�
dB �C �+��^U�a���Z�/k�46f��IJ3pu�Ɩ|;}i���]�^��t,�Z�&�;	o� 6�ܠ���'q���	ނeh�dw+�����L&��m��@�"�o�[zً>��ͩ�0>�C�+n;!?=I�,�Y�y��%L��{K���g@��iN~ Yx��7,�ra=���2ۛ`���+㡟�B�E=����;.�5䰡�j�YDo�|�mxcB�D�8P�B׃�G@-�(��`�X:���=��B&Y ����V���/�y���<�~�,<[��x'�&�B?S��H��f��nvV�a�����W����k�����S(L�[^�^���+t�PyC)�!���r	�w k�P�,��ĝ��R!ǊI(���B��Nl�.��tzpH+�	���-�D`\���b�S��0_�����hk�C{��u��3Pj�r!�9_Ѵ����y��&Y2YS�[�֣b1I�X�a@������k�=��c/��iÁ��a�D�X֮��afn��wW��0�}R"���R7�e]�DTk����ΰ� X�����L,'�Sa��y�A.h%�1zņ����g^������J�N��r (Gىm�<!ϓ&n���5��p�p�>w��ۗ���p=[�j@U<�(�&�p�@"��`�8��՞�#�jD����L�9�Tp_�h�#|o����í�N?�=�L`��!%��(��Y.�?ayD��tpw�gd�ךUr�4ֶO#��\�S�v9G+ �Q���I�h
�����h(���|q�q�g�`���-��E���dw$8���� �W���Z5_ ����e'n��#��jT�7�Z�_��v?D����Fc����.��i�N��X�^��?��P2� q���~K<UeІ,�B�����n��eVX�M�֩W�o�l�xhr:�
<I�Ha��?UT���Y���U��:�U�����ѯ�?ph�bQ��=k�S8�05m-��p��@"�
pV���,�,���3Q��v���k'�w{���H��L��Pw����IK1��<m�E������4��m{iUۙ�{xY�?z�w��aaN8+�LQ�o�1�m��i��_�gx�Ҟ����@?�2��ՃC+��ݯ�y\u{��6pr�����|Й5���� ��z�k��C����H�l�1�!�Y'T[�ӽ�e2[��B�95���ҕ���J�٧2}���H�j��<A������o�"8�Ԑ"Qe������=y������,7��Kڪ��V9B�bW�{vj����቗0H-��B{�M�όrn�S�O����!���\E5�]	� ��>��}��EB��u�ȁZ�A6�%����n��{�;�O���u
dQV����⪪OX�ݴ �m�^h�?��,�^ƘC��S;��{늿H�����>V��Cv�/��Ly�=��z!䋼�.��yQU�̈�N�/����#=y[e^�i��g�����S,qXe�$�+��/XFw�����F|���p��q�f�� m�J�� $�>��E���7���.�`$.5\BU.�5�7�N�lf��rlЁ�P�~�v�'�2z�@/���J]�;�8b ���*N�*�$u����d�vs\N��0��G@,%�]~�g�,���D��_F9й(�gZo0ǈT��e�.Z�t`���Vçkj�r�"�|	��>L�Y#z����VCY��{Q��$�I��(�Ql�vS��a��E4Ût v��.g<G�o����S0�o�bKj�/k�y��2�L��W��(�;����ˢ�	n���#>���fc�A�9A�����_�@���>�����V�+ ��]xWs���4��G,}j+jn�$��Ş�Zˋ��Zt>�/�&�B��x�4ԗ�w1W�8�6�� �]dhu.
�`c\�"q$*�h.�<��Q+^��z��y���r�"��^
�y�L~a�AsڛR"�qF�Y�lM%k��;ɍ��'!C I��%�Ӟ��cZP���
%�f��[��������g��,��t�H�W�o2$3,��Iխ��d���︰���3�	qp]�)�&,����Tm=��Z����k�y�x��L�<3D\|-?���&\��ۏ ��[����y�1E$N�j�8�ϵ:EĽF�%T't��<T�|=,�R� t�i�VO<JUH�i*m�?({ 7O�J�j�|��Eg��)/]t(x�ux\Ǹ��昣^6(�<�I&?�O��o�C��L2͆ABtA�*Pu���`�k��N��ڜ��YM�f���XOxt-tha�����h��Ka�T]5��L���_˲�����bk�+��l���������l4�zU�OϘz��*&]7aó���	TQb�7�DK^l�K۾�R�O�;d�0�T́v���5��(�ckI�����㚒'׿�bs3�{:[͂iOeH4��4
-��C)�����j
�a!�$�^�f�0~%�B���c�j�kI1���9<��>4=�T�$%]YU�J���D��+�re�ƴq�lF��N8��Lp#jS�y��hd�4����K�j$?�,m.kEz!�7�0+?���T31	?���<o!8QkV���u�*�^�RƌրC���ϻP����?��|^�!�+�a�#��2X��z������@��b������3S���ZS�T�	Vi~.��d��L�qN��"�6=s����-_�x���0��Q��ƜQ��q�a��r�˰�J�K;�/[�Jrٿ�|��.sQ ��K�s&f�}�[7�zG��4b����ځ���"��`��҇8%:wV�ٓ��7U$�V�/��a���!2��^`"�Z�D�ɳ�<$�ra��T�c��Zڅ��{�O-'w���Bo��B2��z*l[�p��q���N �:`�G��7�Yd@(L)ج�J\��wA���G8�F��%j-������A
�R�8px����8��[M�V|i�!���E�����.'�yvJ�38V}�4�Q�!���P	ք�M:ʹ���ENn�i���4�1���nKԪ�qT ��7� +�H�BV��Q��g��H长��-@��o�,�S�����\�i�������,؋��8�lՋy���;��؇|�AC�m4�s�,n�꺏*�v��5�jGތcgS�L ���K����l�zo�T�cנ��O�ϵ���%`���ӷ���6����ts��X���p�Ɖ�H�RU�/����)S��"s��ɋ!T���w-J�������хw`��M!��0�����u��������\��-1�o����qؚ4�L����b�u0ș�#Z/��9@9E�3�����6��j�xl � �ा:�ÿ��Y���r�hF�����A�2�l���_RC,�Z�J�h��He�KHv
օ��n�S�!O����#�}IX_��9;޵>�CQ~Q�����|2?-8ǂeC��Odt�􋨋a{A��%us��?F&8K�� Q�:�D�>${ܦ ����yx�n�Z�)�g[s�ɧ��0Q�1����,�2Q������z[[$�5A��T&�f`��Q���\�b��N ��M���G���d�c`">4�"�F��`���{�aT61���C7'uu.;�L��m���z�1�,�w�*|@���t�{���k�GVL1�|o)�9+d��,�դ��_��<p��1w{����b�l9�$��C!�.M�'T��/5�H�Ådd�!�vЀ;Ra�����nW�ޯ��[-֥��a`Pγ]�.�<*X���8(�LQ�P�yOE5hw�޴�bw�M?�F�Ie�V��x+�<����_τ�o��_#ǅ�&0�r�.���s|����c�z�����DV���΁�Z�O����4GO�>?(�Mf̅��b.�zFgb�ng�U�*$,6�>�E��(v�x����.,��-��6�Z�k���$@	���Ut��&������/y�Y���G8��pk�;;�2e�݃б�Fy�e�}�0Ɩ[13H�4�k���ɵ����r�^��~l��4���B$W�"��0�Oo1QzR�	��2�������*����v��?2�Z͕&���,!u�;-*o�ּ����Q2d�X�4�>���@���Lr��Fx3�V���2<NAh�ܞ��sYj�Jӱ���Y��$Hnm*�����?f���7@�� 7���ܢg�I�V��:m���?��in��C��Z�?r	����ZO�U!2�l�q�i����H�\h��	E���d8֌am7S+c^;yӹ_�[.�Ԫ��z�Zw�"�X`�.�K�q<��!Q��!j��J�;_���鶏 \&�8ZՌO�<eL������<>�3I�l"V���R;��Mt��1��Q�hhA�Z:�ʎ�=Qق*��X`wWWÉ���Z�՞�:se�A�(�dTV�f�#/&�嗐S��������:y�5�ι%�1����X���������'A{^{�}#�W���dR@(v���rє�V�5��f�e������'GB��É�& !�&Aq�����u��l +q4!Z��cP��f�p��-Wg�{�=�6�@_�$�+h�qnt\�\�
���;OjZ���.4�om{:P&���U��]�k�N+���>�x��/�
��N�|��GS�� \�<9$����>>���E|�1��t��# �@s��vl��q��	���'ν?n��T�����c6�z�7$y��Zz��w�c�pJou"c���u����o��x�ḌB� V ����$��ٵ�%�i��BԆ�o! r�� �WL#�(���t�K����lU�`!d7�N9VGh�6�ۜ@��-����nv<6�\��-m�D­}13�ԃ �X5�>�]9'�҇J�4�I�W�M�$�z�}��`;���v1�Z ��(����[�X�_�1J������{'P��F"̵�T�Df sZCt�Kh�է�/�`N�)����.�b��I���hjUˣ[:���M���F��US����ۃ�|�����{
20��� c�T:ԁ9{d�X6>ʑ���@ys+�L	N��V	�K5oT���~�S�I%�۴bKj��%��A����_D`��B��س_mX2q����>�|���9=�a�� ��֥T���3�_m�p�����L.�8-����VE%j��:��ҝ�2�dV��L+��M5�5*�}����/�V8/���&>�g۸U�2V\	ƴ��p�Y/o���Љ�L H��G�q! Q�!x�8{{f��n�CPnP=hԌ��40k.)��G=��� �����
\���$�[���B�U�3��<����mUL%ެ$�N�iL�(����@��C��-��HX�o�����M�M���h��J��Ф�X�B)I�uxǘm�h�CĈᅕ��Ȋq�#��/X��a&�U__+�����I�~�˘�Ҧ`jG̑����tD-wLc���Ȕ�VR.o�����ui�yG�jpA��-+" p@<�!�W��l� m���ȿ)ڭ��"Z�6?��	�"�W{���/Ol}Ĵ�	׼Lޞ+jXz� �s�����X�մ3�8g�.��T/�~NM\�;F%��Dg�a*��\Sר�s��x�Ά�Ӝ��+���>�$�!7k�4<�g~¤��=c��|맾�Qo���tV+* ��,�6�w�,m�𬳶²�;U�|��v��]5Rs>S��Ӵ�d��|4�o�>�n�0Yz~�j�<�3�]�hըU^ƈmI���x݉,\�:�ѯ�/��T���L{i�*�I��HdR����fV7tK��O}]�Ǳ&.o�)��ng��?�+����v>?���;�NN��+�\k�}
����,�/^�,U�wU��Mg��	�t"+@pc��A;�CM�'����veS��W�����v����0}�r�9��
���/$R�գj�'Q9Q��W�J"O��_�s��B�D����㵫U}!\4Y���ጦA ��\��G���n���,M��pCX�)-����#kY��	����%�3i��ЧE��Dj ��_9m�EӢ��
!��YY}ګ*"ג޵�i(J�t���b{�O��
������[�-�Q�e�+ʖ}���i��թ�들�{�A6Ղ�89Dt� ���$��y�M��Su��KDi��){=�u�KmԨ�ހ��Tj���\�/�ՍE��H�ii`�0qT{�^��'������BL�in;��悌I���~��+��l-w���'�8=��t'�>��b��A#E���j�L���(�X[��a�d�
$lD�l!�d?v$7*6��|�5���D�&G���\{#���-��~>�Qj��&����fI,�J������Į�롣5�O���m�[aM�D��!� O�+�[x�D���oo��|3�S�9B��s:�۴Q,Κa\�>,���0~'��:ԃ���3��cQP�d�5��P�G�]�J�;�rզ�ݹ�d�-���N�m����T���!P�k"RJ0�0��t��� ��Kz,i�(+Xk[[2�#Y��Ӓ���z����Gͧ�>��̵͊4o��(�.Kbt��ͳc���e�%N�iҀ̳�Ѐ�ϒ�߄��1�˒�g��뤭�C�߼�T���]Ɗ�zg� ���V^�]�Uw�Q�[��f��	�^=M9p
{i��Ű�çZE�������'̟�Z�	P������	�1�1ܨ{��K�"UR�c���G��G63K�¦�l�xd5����̓���p.3��Y5���c�4��v��5�-�Hᭋ\	�+�Zl+�|ѩ���{�u���<� ��� t_N�4c,��Ĕ�$v�-�Ѝ�n���-��@� 4�Fj�s6�/�,ͷ���	��)MWL�tD꯱��fO+	���I�Yk�e�9G
a�q��?��"����f�U`���7*7�B3�#La@������(��lc��۸ʆ�g �?�����$��j'+#�bj����w"��ǉ(]$-܋��9�C��QR��z���rde| 69E��j��m��|�w�&N�&�n�I~04\_�lw:�>��M�C���9�)
��gJqo)@|!U�#K߾r��u
�X�bc��>8��l��
^f/˗_9� }����C*ZۛQŋ�i��8a�+JB��4�,
��Ż>	��m�`V� ���+R��,�
�3��v_�x����z���'. x�6�3L�0Kj�kB�C_�
��� Kμ� �9�|T��h'3��D�M��,Ή�̡��_y2+\�.Au��_X9r�"
<�����Q�ݳۑ�l�5=���!�����3���Y�4	���+�&z�=9�v+��K0��Z!Cj��R�AO���@ثL����7/�����c[��5~��\��J�Y�4��I�̾N�Wh��`�u$��i�������\q�K�Q%���n���5!���E��-ȪI6��@\βקmI�8i�J)��|���uV�-���$%�l}�A����8�����(X�y��-���~����;Y�- ���Uqk�a%�z��˫�斵�ʍ��?������=xKAY�r'.�]���Z��%dAL_���$�Âq����)Q���P�=i`�����aa��3H�E���y���;e���=�=ƈ>o"w��F7<J��(��k��)�ٚ����D6\��5�;�q�oA*e�����(_�����y�}�֏��LK�=�3&���P;�|�me��jt!{��=����q�c�$aR�Q����
bD��>��fd*v���Xb8!���*�;JtW^���Ayp�rC;$�拈�X���香m�����4�_"c}7���ư߶�cʆ�4.��Ð��y�JIm:=�%1@ELWH3�8�9S��hY�T���O��}u]�S0K��nt(�$x�K8��h�2�&��
tl+�xae><��;>�nV�}���<rA*������mGg?�B�5�8��*S�D:����7"�H�l��W���5��U�����s=�C��8�d��s�l��DJ�	��}İ�UO�#�*���j6!����%�-�8t{0�}�m�1�Ry�f/"����ݗ�O��K��N{�	�B�u!�I�H�yXa>�ܯ��oA\����b����7� �0���B�_��������RC���{�pw)����o��:{����Lgn; �
�d�)f�XTƛ��/����~���F*评bł�-�M@R3`q⮘�YB�.��|�}��\l>A;5U<5��;��G�pծg������юg¯�w��*�+��(�cM��0�Ĵ��+<�̬��ݟ#�����W��"��s��'K����}fS	��]�O#�^�)��6[�$ָs�(U���E�f�poi.]3e�"����cQ��(H�����4u��#��4��t���-K,��}��l�;//�z-&��i��T|��;+�{%j04,AÌZ�Cۏ��וȉ�E�X�x�XH�,w\�.y~D�]!��n�ْ@E?oUƟ濶{����9�4ں�[��=�EV���}0��o:3$����,�N��)]a�Ա� �}Y�m���ܴ"KA �.;$��C24�؎��ܨ�%ұ�u)��a��?5�]8V!�"Uڮ�'�a!4m t�۹�n� .3�>>u	��]��MKU|��/�d1��ZF�w&�+\�f��46�;4<�L��׊��FlI�p����MO�/�7I�-]M
����V�K6C��9�n7:Y�.џ��4�誱�U����.tѬ�W�&����/f�=/�Ą3�ie�
X��x
.��E���GFQ�����ȑ�ݦ�*I�?%�T�Q�}Cp|�,�����.D�/�� wDݓ�3�Z�+�����/Z/k�;���mMj��$�X��bwf�uYN$S�b�KL&���	=�����N��K���=��H��3���N@��39�a��I������Zs����a�i�m�אU�M�*�;n|��ǆ.I(h�)]� �8~��������
�I�H>��8����07�����i��U��,h�D�R���]cd�R��J=�	����^y��}�|4SIrU�ȨI+��Qo\ �L`ժ������"��/]��'�C�����ʇ�Zk+,�]������s��p{�_���y��^�7���`���ԋ���C�?�>��[�;�8�������w!��9$�u5}~��>iG�5��$���l��;&��۳�9a���D����t��U�v?���\`���/�����l�'��I���K3�"T���C�Qt}��S��>H>��J���+;l�&|�=�?Z6���3�Ƹ%CHn~��h���fF�v�b�$���\�4�98�Au�܅�����"X�ث��	B�)���.Xg���$YO5�u�'D����b+�Gp���7YOl�!o�}�ԫ��u�J(��6-��m�^|����)��;�R寮��ʹ\��d���w_��
�䜭����Rq>(�-MBp��}���ks�������*=��*��.߀Xʥ�|-�1<�TD�34�V�ʊv���?�W��%_K��"R�g������Fea�~ �Q��n�n���Y�*�#�-��J,���6�DԦ.��b;V�Ws���_�w�rhԶ
G55�6��E�a3Q�o���s�loe�$�s�j�Ʈ��}����7�h�I<~���9��Y�G����7��vd)E+�$�ǵq�ŵ{� �t_"S�b1�mP��Nq>���b�N����WPeU�r��%�F,�A>�9b4^��,Pbӝ3�b��#�$9'��t�{�5��Su/�J�q\e���'���Qȗ���ב̛���~|s����T.� #��� ����I�i�s�s��)��6l��>d��!����)L�f����x%ڡk��C�:��BO�?땏�Wm����ڐa��;ѻ�,q���y�L��ލ�Ut�1�%��˼�*XT����U�����n3U��$�V.��s���ґ�TBc JLF�Ջ�?"o��*ٶ�$}`��e�|p쭈@�8�����h������$5�2lrWT��y]�4�Ζ��E$T[ԗ>����i���t�0���<�Q/�6�{p�	8�]I��6����0��T&�8�8aV`��.:1]_V�~N���C|������`�Ci�l՚�د�m!z"�L��j�B3�Ï���� �4��:P����L��#���'0�4�P�lm$���+{P%���[~<�O��Х�j5����(��+tT�$�D�<�\���[@s}�%��n�n>!|)S�����PQ���i���]�l3��^�D�X5��\A�ֶτ���3��?����К������@��O���yi�&�(#��Gx�oe4��&��|�܁����e-��+j(@d��ku-b�H6���Ň�S�x2C�=P��i�(�}�N�b�2ӊk�:}�9z�'��Q�Ҭ����r��:_���<�J����MW:�k@����{(wN�1*��)���;�N�d�_�ܵ�	��4�g@I�?�~��KpdY��wxJ<!h3t��yi����J�f��,&��\ _b>�-�� (h8~�[w�v8F��ݵ��HȞ�0�����O�đ��w'��iL�O�-Z�%�,��d� C�#�F>���aq!?ʵ� &9�o���c��yv�E��.wY �㻖�&/D�Y\�$���F�y�rH��l��l�������#Y��4G�i���)�����s��Ȁ�s��wz20��)3�Z����mm�/���w�tSKRxV}� qi��|��Z,�F�����ί��BÒ��M��Z�W��cJ���G�k���ފ�bo��|�:+X��[�1������*^N��%H���Xd>�OL����-c�a���R5m�?���%S�Wͼd�2`�9� Z� �X���*�P��<�����֘�=_^%L����rʈJ4ʓ���;��/�Y��0x��H�ɸ-�#�6�7��.�6�6+f$r��5�Le�'��h6�3N,2�V�e�b���Y"LK��^�o��2�#%��I>O%M	�ﾈ/�g��U	XXu�@����[�&G
��TӑзL_+�U����Ne�w��j�"1D��E� E�K���#�^yd��w)R4��>cS���MD���Ҵ�$z�k�dj�H�>r��za�Ig^�'(~����;[@K���&��z�[YŠ����C�*�1}��G������<HK!��]�Js5
����8����Κ$�*�_i�%�E`�XN�?��3�9��>�
����/�k]�i�ű����iq���oϯiq���A���&�iyM�l��e')��/b��>]^`�[F�'C�Zp�hZ����c� �~�(�
Є!o�r�Bo�������ƓE{.��61���&Ayjӥ^Ʋ�OAT�!ǡ�-�����t+4����c�z�7gH�3Î
��Q�>�0,?"г~kaL����
�Dl�|V�\L�>��к
[a����I8K� @�!��c����)����j�F*Ȟ�>�j��C�*���	��ʑ���N��(�۪�^g:@P���i]Lp�I	�C���(,�d�{̥ƍ�O��,�K"d�P�	v�o�/������I�����[��7O�2�p�]��w��ffc;:����P&O EtΗw|ؙ�ݩ��4DF��&�9��qb��S�=s0�4E�2�EQ�&W����X�K���#4�[gO�p�E8�Չ��dM�@�,�y��Y.��E�AP���J��>jC�n�(�p�SՒ�b����p�$����Y]�%��o�z�Q%��xu���3Xs�����R���W`����#��ι����xp�a�#������΃�����n@� uk�v��.����0���R6Z��3�A ���9�����BGWUHm^�넲����Nb��a����]���8)��"�<�5����C/P@Dw��25��*n�y�c�n�R��(W0��wZ����<D~�r���*Y/�{���#]<1�2�� jD�YyFYfV�xϚ�� �u5m�%д30n*2W+�͑�)b�Ʋc؛gJ�u����M�oAO�(O.s�(�*NR��N���ݯIk|GxKh$�^��&�<�2a��Q�a�0�;	�%Q�eKгW��#G�k�VխҞ	�Ld���W�3�7������ڝ�k�i����}]Q׭�h
r�
E��Qb���%c׽"c��I�LO
J��yzq�����`y�C�	���HI����Sx����׃��>X�e���	�7.�����)g���֕�Ķ�'���f(�"�b��w�ׁ��M��T?L^RZ}d��i&�$�S� �`�����1V$�B`jAǸ����Gq�c��n"��\;[��G��J�yI�8!��b��e�oo�&�Y���˸=V��\�Of��%�s4�pN�e,�5=iBC#���As��Pk�?��Gj��9�2��v���x��) �x���Ե��N�a��)�;3�@���n�a��(L�H�S�VQ���h!a/D>1�!���ߎ'h�*xK\����C�43r�:�u��"`7E�=�!E�⢴@r��� �J����|#�G��ή`�L�#��"�:˭3�z����K���%��$���
Z����8��|Ôg���=\�1��I�� M�!���7��ٽp����b}�G
[�TB�9�$�6�pS�ߧ
����ֺMa\�k�u�lzx��֜%-.I��M!����V+�"Ȃ���9 j�rO�q��Ca:�5y�����5�kdd�T'Z�tOA�Ԍ;�P����\����Ýj�W�o���#5�p�aZ2�5tw̗^n�%���u�����YV���G�k�)�#�-���	S���EK���&�5n�}� ��$a�J.)�0����Pi]Ufe���y��2x��6�:��р]#�0U����T�������A��wa����Ӳ��{��25ɲ
(����?�����W.a�C��ߍ�}�E+T���y���۩a2VB`���#N���"�G�����ob�1��}ȓ&sR'0�7g�������?����=
0U���6�����/��z���� ��^,��D��bt 08s�$ŝx��VB��&�:�I��ɜ�O�#�߭%Fs_K>�	E.�zeA��8�Y��|@���Ut�~�� �"K�_%qH>��������_K��U�S� p���X`z��>x�D����'��/˻��D�I�e�]��ξf�O��2.�ZG���s��ҍ�_��_� ;�nA+�ަC�`� <���NX�ԁA)�Lg����x�/|>!/t��ؖ�q�v۲j/�?8��䣯p��jOV��1~<����c�{��U~8�Y��=��
�,�l�I-W�p����7�E�5!O0p��$�b����B�V�C�UA�,�H������2��� _+ر�vs�'8#��#�zY��}�Z�.��b++^eʥ�[���x�����}�~�o��\����h�3{���B�<��3l���T���/��&�"?q
�R߁+B;�}Tk���dI[�2Z��m[�[�]%ү2�#�,ӈ�+t��V���6�5��3��3��|J�&��-��"~��a�ĢC���t��i&����.3YєiIXR�����s}LV8��33Щ��=�c��&��Ut����u܃3��O����it���l�P��K=���l��\���W�9��,�廊�t$���&��8�'끾�<j�ZL�:w����Iz,.d.����o�4#�Tǒ��q/��ai4�T�\懥0�dX���XɊ.'D�?3��7�}��� #S�V�2+ ��i(�՛j�<�$�2�HV����	>;��2�W���m�^&� �k��h߸v~GY��^�o "�,x���g�k��|V s�Lx	�X4I�Ʊ����<����װQ�7 ��^��j��|��s�\�,����¤�fk��:���ךp�<����6,K���z�/�e��<��EF�������Aև��>mX|*l{��2��Y��l���|��8�,�jV;^����}����	����r��zȡ�ۓ��N�׼ƈ.�*��{P�h��E^-}��P�, ��s1���s����d^R���L|�J.B���`*j;�"[ʿL-gl�~�$�?��X�@�Α\�F��Aa���L=�����Ӑ��?����!�i~9�,o�RʒƢ:�����^�0�c����kՖa����4��@~ɷ|/��)>XA� _@1���+l�N�����V�ΥM�T�q�M0궭� Q�Ğ$F����sp����~��������>6ݭ�"��:H��cg@x#�i�S���
o��%�=�}��5R���=��=��.{�+�JL}����>�� Ǫ���Z�ԙ��X��"�[�����x�_��HK�L��h�w���*�?n2�4�����m���R�°%����$6�в�F	J����B������ R̤Z�Zǟ2�@��ؿ"��M5�*�� 	-��<{��>��g��i	��}1�C�<�DJsE[(?I��/����5�$'���~��z�ω7�pX؎"P�� ���s��P����u⿮ٗ��~ڗӳPb�#U���i�XκR"�D�t�=���c�3{k�u0wӞ���{777d������#��� ¦�8��I�B�d62�(�7W�ruT�C�U��CV0��:q�ű�а/�V����a fJu�f�[�P�"7�-4~���ғ*]��uLsHP9Q(z{(�|)�1:R$G��}K����-������}_E��t�GAѺ��!�e��E���Y��:! ��¥����'AZµ��ZA���W�Q�{2��7���z��PʕP�� b�)7�ݤ��b�آ	  uE4�a���v���D6���!���N���{�Z3쒆
(�/"���o��M�~�1fY_��BD�L5F���F�i����3�wZ�,|��!1�� 4֚�S~`!�%5�	W�����i�8�Ī|����96��0'H�p�A�^���y�I�B{��ۚ,j�g��"R?����䮮��I���%y�U����_�d# 5 y��\��sU�O�ξ�;@� ���')=���/W�A���eh�a�J�Gi��3��n�z��W������w.`HȲu'��{%֛�+�ۼ�"'���@�n�,���G�b�<4�P���a󻀍���&�N��*?yt� I��z��(1�G!*�)�|�v�*�`Ϯ��'��.�g���p��S>�w��@��P����&��{?9�J7�w�ݸ����h:haI�| ����hh���<7/熲�:�Qū\1�����������^����n�$�����R<]r�?zb�_�;�)�M]�(�d���v�@;��}�<k������X\y92�m����|h����ʺS ��r��+���}ZR��)�?@��58��~�H����2\�d��9~[��pX�+f�H�k�e��@�y�Y/��������n 9�56���̉���Y?�?���>Wd� �X�W�Y�\���d�~��|���?^�~>ӏ���F]�S��)�	�sO��]@mT��ߘ�I��_Y.��o)�8B�ʟ�fJ�$�|����o�2Ns�X���^HHЈ���2�Ƭ����I�G��Ye�6��� �J�<;D�D�xH�Z����Z��?#��IDV&�Y�\`?4��ڌoK� >�㎄�RE�1a�j��5�(顱�a3��UnLu�T80|���*��D�{�Mt�N&�U���MSk�fu�;�}��}?��Y�#cU���S�\d����p�|ٌJ��Ji�[:�����A����r�]��&��d4����n����l3��H��$�w�������6Y��ү��|~��Z�!����;��^TN_��^������v;֜�j��=I�����J�_}U��A9"A5��8�^��a�s>�'>�ɾ�3M���@��>o)c���k!h�����"����G}�[�M}{��e����k���5��7R�]'/�Q	Ľ�Pn�"�ZR��sxP����9DK���=f@�� ����K�'*�q?-�%��Ag '�>�z�@��,ľ��T�ޥT�m�E���DGK��x!,8���YV����8���Qꫀ�����Y�t3���N��E�㓊�tWg����[ Ш�=W��i*Na� �g����䏀���h~;E�d��P��Gح�ӆ��[wZ-�k&��s�k�/61�X��XJ�K8�Wgq%H�rx!U�F�\��c�M<cfN	?���yLj-�!��D�;6����ޅ��]�c��F��p��g�|��tn�E�ڿyr����+�=��u���:���T����@��0�w�8�5�I�� ��\���S��D�e�ʿ�������Y���1r���.Oz��B'����Â�(�����п+�ڳ5Q���@��]�&��˴��> Ҋ��S��@��T�Z����í��d�klنA�ir���D"�W؀S8���G�b����Ѡi,:��;�M1˔:����:�#���}�/(Fwml �c#^�y+l�f@��}�>��rQ{_�E�U|�_X�0�.�������UѦ�u�3�[���{��Ap��tn)��b�;��8h�q�]t���?��Yu�_ݛ���M�Μ��%K8�����:K����h���- &Ao����8[����g����a<,��F��)��ëv�0�ۧ�x���AWk��cJh�4p���D��Nax���*r��������z��x/��V4��J�k� n?0�\�R�:>�g���(GrB��gER��^-嵴��W�aNЄ�S=���c�Y�"[H�!��Y�'_����ϐX��Zb���:T��8�\T�jp��1D5]Wt"C���E �E;�f���y�7e���N����"����Ϯo�-�t�x�2w퍗�9a�{1\e��2?��a?r	�&��	�|?qV���ou��OA3�_:�!�U��j�+�!F��~KV����wIǻ�ť��S*��BY�qUiJ=��vF�����Uo� YcP��̽KkȒ��y��d^�πO�aym�+E85+�:�c��4M''F�`.��'�j��q��ߐo6Ȃ��GS[du�M\!|S�l�8���^��&h6��nΖdI�nո-&�9Ӟy��*�PƆë�X[���y��J������uq��BI��b��TIEUHJ�/S��H�+V��@�.�M�'�*�.��-"QOO>�:���U�7�tӊ���tZ���������"@Blo��PpLb���Q��d� �������[�p��'�7�$�*�S�!��)pʳ�n�jR@3V魎��Ͼ���p�5|<s��|�bb��f�0�!B���nr����r���|,.�s��$��'�IsNɳ�Ny��C�y)��L��b��W��K�m�x1�H�²��-d��Y���}:�(�*�R�H�}e֪��k��z���S&ۛ�I�����د�2�!�������}�p,����{�z����޿�}T��lP2Y��U0?fTA@N"I[c\��xմ�j����J�\�b��N�<f�涖�ɂR�7�� b��:e�]ǹ����ƌ�@�s��ĻP�~���
wF�N�g8�5�;�@b����=��S%�Ht�$����K��+}<ը��-��`7�vA$����`��J�.~Bm#�� ��׊1H�h�q����w��^{��E�~�=�%��qI�9�[���;�>ᩞݞ�8h,¾"u��=K\���(xDv(����P
��/���8",�q\q�ʞ�����V�Fr�y��.UW�:(|C8�-Y!Q����q�~�?�i�;\������m�R�nd<a8�;B��J��ȦI喇��8�*�LP�y�R4���'�>7��D鎂�$Cb���qadc�Y�0��%��6�(I%\dBgV0^���[���^"o��g�X��>.�	˪M<	sRǝx��J��	�Ƹf�He��@�B�yaӣX%M�e�Ճw-ɦ��T�Xf5w*� +�O7�.�v��ת�A:���V�@NG������pݻB����c�E؎CI-aߝ��7�ݠ��+e��ײҙ9P1�U��ja�(4?q>��*9mL��Ha�aE&� ���o��{��?@-*�{Ri��LR�_�8+[E^�E�[� .�u:�(G	S�q��+e�	?�����������鷙!�}��?�2�G�B����r㧜���}{g�RE��7��t�ܹ%��Õ��$�=(z�?����*/�jS�����i��Nx���]6p��Y�?r�}���N��!iq���5��FY>5]����=��G3����a�l0DSH�����(���nenu�5OEa��L;�0z���Qv��ƔN���?Q�x���{�K۪����PC��x0�����ېa�R�A�^~9�����Τ�����ˍ&!�Ŭ		���\ �	3C�ˁ}p76�$@����yET}��Z�M	-)Ȗ�0�i��v8��3,�y�"��w� �Z�5���*���"WPohgɶ�� �@.qQ��S�T1��|��^q�Xv�o8�\u�>��������/����[˻cmF��Uu�LӽC������64���0I�8�� �BL�t⺔�2�sD	��\���SjQG�c�b#�&u�5�����N�i��f<�t���.��#���8)C	v�mȈ�s�ܓ�Ƒ�~�����g�G"^�đ�ړ��ĘD��B�M]�Z��ր���Q��2s�B����2[����Um���Y�4�24�|@��-�},�t�x;F��I|�;o�/��qs��&ĥܺ�Gx�6�2��`������'�"��S�wmj<B������P�R����a)��i�(�����k��5�֙?�T���8'�پ͸ۿNH����O���ӻ�Z�z���W�{�w>�S���B���s�=.�����Q��W�8�p�<=RB]ۡ���ޥ�ö�6��ٙo������Ĉ�=Z� s�_�t�;�5R$�06+�����>�p=6�s�bR��L��>01�y��-t��fo������,�T��y��>?��[���*✽�#"��^�]�ks5z�U�yrp�*뙈��xC�^��|RQc�^�3u��.�C���XOh���"���h���4��cc�ㅛMJ�C�C�Ƕ��@�J]������������쩖��0�� �=���n��̒��{��фǿ�n�����J}�#g��D�l�6(��6��|ri�6�y��hGJN��XL��.���|</����˲<���˱�4Bhe�f�B��),��',n�5W�-<�$�m�7Y�f�/�0�?X`�(B[ Y
����^[��PȆ70 �U�6���Z��)�V�$��3���Z�.������T�-�����T-�0��ċ���Ţ�?H
s��:�s�
v����*�Z�>�G��U5�%�z����WE�
;�О2�~�~��t��i�0Me�;�_�R4g63Z�갳l��QÜ����+����x��E�#Yg��i���k�a�.�K��.=�֕lH�{���/H1��ଐb{�"ƙ����T���D$v�#̲D��aJe�f�>���>xȆ����F� ң�m��+?$���@v���A�ZV�m�����T��v���¦.R��	�!���q��
�Í�Ld���8�N�xGe�@]�ZO�~e5������N� �u�_��êto��A�p�Qu��F�ȧMH�aEg�Q�UI��y?U7����b_I{}1E��$�����!a���`�i��o\uzt����e�F^+\��a))U�:r��;�_�4�H�z!��ǳ3_���gF��Exa5�R򐸈���%��Y�]*@���5�Vqr�2*�@| �i��P=�\�Yڻ*'`��*��>އ�x3d��]A�����o&q�����E�h�q�p�]��$��W|ͯt+ҹ��xȗ���
S�<�-Υp9���:!��J�!OU��F�P���ȝ��}{)NH��j��,q÷�:��i����^����ٕs�J�����W-
��{����,7�_M�,+�/cw7���#|�&�N��?�m�-�5�me���jf���^��|�BWa�^Jh�V��
�1�x+p&ѣ�/���e7d-$��۪:�U�HtY/1&"�qf��H����`�S՘̅�%�[��L_���'�BXM��j����)���T�7��'8�^I�1���n�zRma�������2���95�xF
p﵆(|�ŖW��l��b�W�M
^�1���BH1!�s�;�}6�b	Z]nm(5ٮI�z	͗�-�_��y ^+��?���`��O쁝�G{CJO�@@s{f��?Z�W�M��Oc�Y3�+*�b/Yb��Cӛ�m�;���#�E^����ZSï��{���ƗE����ȃ�Uq4��q8�@�C���A����8��.�e}}���ۼ���ʜ���ۍ���H�b8����׷QŎ��ɷ�o�T������<��;�K�l��c���CNK*8^`���0"AOX�6s�����oZr��F���r��Y��ʭ �#@�Y�%W'� �
�s��3���fr��ʖ�.�B!@���t;�?'�\M.�+:�K�B��Ѩ��.\%5^�����I�h�e�7T�6pZ(��@S���`�q�T�oq&��*����[l:y'#Mr$���{�f[^B��;�B ���4纾Zgh�������\I���Og����ժ��~�_�ۨ��������y~���jB�d��φ���Ӻ��͖^#��	�O\�̊�$����/l�/�x����G����[ҵP��ஜ��L���x՝�YP��ʨ��_d����p*�y����z�ό�GvE/�W-umM������yp�3��nj��D���~����-��1k��t�Lⴛ�ٱ��I��hΔ�j�
�8GF��H�-6��wb���=K}��M�i�����֌[���眪�]%��p��gLm=�d���+��!~��l_���lxz��tfZVSZ.J�ʿ��/�"�Dd�w�II_ґ�w�m6'UOoz*������������ƾ���O7רTb��~���a2��_��t��� �?����3)�Q5�(�;Y�0N5���8�S�،����_�\�������C�W��D�
�4�4��c
��k�w�"{%��_���1������i ��A����g�gA��v{!��0�!7h����j�z��>���De}s�1�W���X��S�\�e���u�>��932�n~�
�JQ����]R�.�&͡�ߖ� /�N���(�uOB�0?���2	*��
G�&?�������E�ٝ�ś�nf� v夅�"�B`V|D��9&�܆����0{�JVv_e7�j�K>1"R��W|�ڽ�������%��Ա�6�%�x�_���	��I`�"�mn\���g��`@�r �E�����d������*�� ��&|(u��)���eL�gm�`�Kc�;�/�U��s�T��~ٍ.�\�I�3�D	%(U�d��U��;����&R�֏?uw���D�k��%�qi�S�v F��*�R�3��_�D�u6}������a�51�H6���9��[��	�t�?�ll�ԉ�_�	[�j/a����l��5׊fn�.�� �^c|�O��WO]�lY=�#So�M�1G�6i�h
-)G;.m#�;cK��}b�j��3We����҈��������.`�A�[Dy.?��@�����9�ڪI+)�/�]=`���f����X�LUuo�<m&\Ĵ����_<��(�����E[�	ƙ�4�P\m|��.f-���E�:��f������j=e���C:w����:���]xIJ*����('=8a�?�Vj	ՆN��ʟ�:Ũ�?m+4o��/�S�!���m�v�I4��Nvz&-��)C���%����%����07���t��$�2����6(۴@�P>ڟi�w�V� �����ݪ������Na��Q>kd�e��]���j�*;~4|K������QZa5#�{8hAEX8���B���R�~�n/�j2�S�&@�ʌ���%K����r�6%��b��5�WNR�FU�(�� L���f�;�]��2���{�5,�+*�f��d@�hb~ ���SB��Y2Ї7��g����|�emC���<V�y2<8�c���v抷�:�
 (<�)y��9?�!�l�*�W��Y�$u��W0i�6�2�˅��
�D_���L��e�����p�=�k�j�jm�~<�ʹ<ׇ��Q=����EL�Q�~|�.�z#��������K�6�H�sH���6{���Y�%	����?ib��0;lw�q�흄���ˋ��f=��W���oA�)��������ޞ����a��5���+��:r"���P��wa�f�_�9'����=VD7�:��am�ݏ�$�k�<�]�����a�\9� E����8+�L��s{
�&
�?d����)ӯA���2^cY��c�+/3��PJ��=�g�iļw�46�BwJ�ȉ�3�PC�?�ھ���Ւw���)J;�t�^ `�ꓒem��ڟ��������v�CŰu���VF�k���'�o�,�P�w��<C.�hoN�")�J��̳��d�=H|� ��h��V�|��i�PU�"�/��Z_E�ll�B�pF3���d��wK�t��!̄�-J���LZ��AQ����>�s���<�<�f[1��@>�]�9P,�|�@Ra�2�@�O�����f�?��H2�8�u����F�-#��z
�>��6{��I�������6sl��M��L�M�d=\d��L���6]���M�E�������PR���;w�6I�o�����c(	��R.J7N�Y���\����<�W_�q\���K��L���v�����e���0�� 2�d)d2"���` W:݁�P�-�R;��җ�l{��w�[*F���!걽��?����H���*�U勑��j�.�a��VQ���_��*(�+��R�y�S%j�Ff��#
1��
Fڞ<��͈RoB4Q�ud�>�G*�m�'&�;3I��H�h^�g�G�����j���[�{��^���+B�fE<>�u��Ȥ(g�h����J�S'3�?RL�2���@ƾzd��s��<����g!��X��g�������9u\���a��ѱ��(��h��4�K9=/4$֡Jʚ�ǂ��
�ע�����sh�6ٶ%sVm�AQ8AV͆�����B^�U |1i�yL���@^yG����X1�G�薟�=azL�>7��t1�D&/w��~VL�M㚂ʚ����<�*�J����D�e$��ᔥ$�ݦ�UP�zR��v����0��D%ߡ"]�	��1����v�]M��O^�����g6�8-��;�F/W��4W��D���f=;+��C?���8ȓ͔���Eؾ_mF�2�M�qgy*ѓ��Un��A�u:	!�V��xK(��W�0��Q����ϔ�����!��s��n	��dme���S��B�sD���-򟟨�[hP�ǜ��(��}�#n�V-��q['�Lg��Q�p�V��<x���o��!���M���1f�4�#哖�,K�H����@����1�k
vޟ^f���H���=������]}S���;1��Im�]��4 �5���+�U��Զ����5�%�lw"�����4~+���u��*��4��-V�@G6[딻ӫ��5-�6>S��!�����˟����+G\�Fb�Q]�����^��s	���؟�&ȅ`Q�������ִ1D-� *w�m�8�ϯb�6K:�1;>�u�Z<����Z~I��CQ���d�v��ɩժy���S���%^=��WW"<�~h��,��:-`�e��5��l��@=�ARo���Vn�@�o$Ut����KaX�>JEi2�{e�t/����d����.�t�W���Sm�W��H�l��R>����&9�{篼l�!U#�
����%��
��J|�h�y����+p���^�5	o�_"�Wz<A��2��@�&_	(��������=�D�/p[nY�o��T�����콝%o��,�C��S�������[�-A;-/w � ��'�o%^n�܂O��G��s����B��(��=6��ft�~ /��:��5��y��a��V��t���.ʌ?�4�4���GI`��.3�:+��������ٻ������1A�';����;R�k�ni��*�������D\�.O_
İ1���q��#yG/=���4�㹚��Z�����
����L�__��1:t�@�3��=�٨�����#�U�5���sH����s�Fg���C�T%(�
�ap�p���q�˝���O�������B�>
�x#p��y*�4Z��L(�#�v��g�;m��i�SF���X��;'�$p�*�l�4��i]�y�X�n��ɱ���\�Hȑ�x+�b��~a�����1_R �� T�cr��2O۶�G1g�7���2�_ғ���_зP�x5�I�+�IJ�����I�c���%�Rѷ/��\��JK0&�p�3�=��/���B�w��s��� �%YìY5��x�F�:5�����_i����Ǣ�?*��1+#��/��k:IZG��z& iVjX�b��C�d]�M�3���)�K�����|��.�(��k,l��n%�)+�w�'C?��T[ѓ����Z*ӣG)n�˗�7�})H�J/|Vѱ��m&F��;��P��gj����~���l�X��n���9�Ȅ��hw
8�^�+�C�`����=���o86��@$D�YvC���鋰A���@%��r��^(��8���6� ]�>���mݳ*���s�`G?coBl\�.� ��zB�5ȸc��}.Wn�ȭ&cz�\D����
��y�`��O��)􀇖�)��5�4���
�._��ᵈ�ݵF��������4�NiB1x����(o*|�z�S5T�֖	N�G��}`^hT��)F�^c�x!t�.wq�0�ʧ�+�!�I���,�.����>=Nĉ�ȭ#�1+"X��q(eFR�s���<:�T�ݪ���>�����	���R^�]�%xpŠ�����"�����ߤ ٤���ۺZ0]ŎqrKX_( ���\�{�Un�`�y�oeQ⒨hT�֒K9�2�O&0����6���q�6I �6��,�gÎ���T|����=��H����-gs����0{��7x��07(�@&�8����V��GaXz��D��y�o�J�V�#�e5r)՞P�c���\��g��U��a�2�����7{mE��%{�o:�:��<�B�/�i��/��dȳ9ET���f3��]���:� Ʉ����.����*��n8�Aht���{����M��߿�qu%����wA�	:;h��������K29�m������(3�q�F�q��A���%­#,]5��s!���@��!ٷ7؟���/�9��@��x�gW}�bA
`ɶ<˥?Ĉv(��x�Mp��	�x^��CƩ�z��gB����e�ajU|���ٍf&��e ���_4}�Z�ͼ���.�Z�[� ũ3�OmZم�]���q�j��������AZT):���s�-!v[���in
�DF�%����_���$cM"����k�~/:����8<޸\�N����?gU���N����2+D��jE��V��M5caa��r$�=�9M�<y30@5�������#���z��-,C�3�F@I#��h����f��w���F�[�Z��6�k�܅@ˆ���i&y����fS��WxlO�0�/�����6?;�*��z
u��8�R����df�{CE��q#�\�YkN��k>:�\�~�;PmڰB��2���D���0�T/`�ow�z�#�;N<��/rῒ����8SM m��T��l����K!n�V�G"�7(�Gz7�c���|@��e��G��D�׹!O�r,�?8��.�M������.KUA�k@�E��G.���"z헧��f���O.�`N�/����_J�:�Er�XjZq�1�|i���V�+�8�Ϭy*��ϕܧu��-W)�}��SF��R#ͼ�����,�����<�G�3ڽ��=�K�w��r���]G�##!�x=��Yn�� �/}:F�r�h-�R*�U���i?�	%����q��#;�ƭ|u�WP	e��N�#;�ߜ%j'���Օ�_ӌ��)Ν�4g����{|s#]��2�l���-�:*�p���	;R�r3	�jT�`;����^O��g��	{�O�lO�)��-CwH���9���0Zz�Vt�����nM*��S��T���;���]@��0�VJ��gj���%�8�8546h�O͕�O�_=�FG� C�C�
�ɖ�+g����:k�5��T5Gu��OP@�r��������Z���r�������a���V�T�M�T^�=�q�� ��r/�;h0�x�������jG�������*�n�$W�1�������ƪ�/9�� �(T�ҁ�s�=��7�CD�1
L��"�zG�.�A��z���А��s�;�é�uo��2��#l�q�&�U�%��!���xR��aw��`͐hyy84���:h�&2�L��w6C��������V�LF3h-�l�2&Wf}���*�_	|��|�-��{�9�p*����؎��4��c�.��J�g�6�J��b˺��K������U�L�W��쾢k�� @n����ke���D)�FZJ#ӵ>�w�7��߀5sa��t���6��)��\�4�%�{��V	$}��q��?eU�3;,Oj�f�����2�%�a�{�be�����V0qj�S�T���V��2�<ߴ�i�-��}ͬyV��;��uit8�x�<�[��5�8�E�Z�6I��e��!9
�_�e^���ʤ�CY�G�r�a��WU���'�1Z%�}�W�����p@n)��P��.���BD#2�U�����&�{&���և��������%�����s��+Ow������T�{�h1��c(�1"������.c+����Ċn����F~P
�c������R��f��,���Ԙ9(�X.�e� �t�ځO�p�1��UJ�;�Sy<LRZ@6%�A�{.��J�ҙAs�����B��L��F���q�� ���(��K��,���֖]M �c��Xem�|t�hN�ĒS��a��c�}h+����1G1�2�N%J�!2o��1%�;�v])�=mε-d_�*_�v�k(	��#s˂)n�X�ܽ�{4����1j���s�<+t����� `v4N��s�/��Kv����x�LI�@����`�_��8D.GK���_�߰н_���:d�#y�~H�(��W�xުy:�x�t �K\�]��G=�N�'�$�UHP�A!���=�����#�B���v'���)j�N8��#2H�5���z�N��f���a���Œ��)�w��T��ٴL�fo��'
���T���`��E�#� ��K8t��,p�$�!!����C�Cm>�$/�ko��dZ���5�y��h͂�3<�q ZP��_*/���U7�O��D��MA�
7���'
��)xUPL�`��ȹ�'�|q�?� Rt#9���c�0��i�K�3��4ҭL�n#õ�C_oA����2#�I��u|v���w�sc�������F-��Q�*���a�L�T@9MlY4�>g�zї��PC����I�l3�1�������S�c$���@]x�oB��R�3ûFQ�Nj�;Zl0�/dJ��	z���R9Cdw�9��[b���^�7�a=\�զ��C�KL��s<�L���R*�K�T��2�qlQýio�W����b�Zs�Xs�m�9J��r�T�Y�2^]��i�X��K'���@���/��Uڄ=خ��Ń���vW��Wj7�?2�Z�qg&#ޯy%�����|g$+��@�P+2bp�8ĥ��$&�\������O�U��b�yg�_� 9�}F�ٸHP�G��W|x���a��8�Qp-�,��7�����V��l�0���+���D�Z���6�����`�ǽi>F>5�k!�~���Pk[�z�� �ZDQX�R�����g��
zc��x��,>,�Y��%h'��ͣ��3�7-�]�r_)aF̅DL������7A(F)�]�u�`}?�WB%��<�ɹ6�P�����<h&�1�^sY�~ ��"V\Л�C�\�m^�9*���1w��G�ܞ�m���~�
��3��@��~��`��HF��R	�*f��X�q9�n���")ʓ0R��Z����h�]����-�>����a�pQ��bA*�.h�cݑR����:��N�?��|م%��voF5yS��뿡����f�>/����s�V�@�~���Ghay�/,
�J�<g��+L=��bO-.�{ù��DV	�'�4�n8~��'���\�د���^�4�Zz�P��c���7*V%��?��=�m--Q�m���6����&P	)}/�V"�{Y i0O�f�ǧm�Acsy
Ou�&`m�[�za*�U���|~����&<�� ���?�Յeu��m;�^C%Sk��3��`Du�%�<C���i���]�%_Ѳ\T�Й�lk?q����w�j���WU��t���!A�<F��[z}������8�E�8�R��x�� $� b��px�z�� ?���ky�� ,� s*Ǯ+w1�JE�gR�����M���r4��[`��N_��Zx���g�'�q�q0�U`?�g�\�;$G��*�Ȳׄu=����wy��/D-�Z5��m*q�jh�����_�bN�����;rsiG)8�]���sj��9��W�0�l����M�N4 L�.lY��$B]Fwʖ=3C�n��:�O�.3�P�&=�O���u$���Ђ�H$(/J��A�:���aBd�^;!�c�c�3�p�zA�U m���ޠ:���]o�hT�\ʑ
�����!>'r՛.c��lr�
����q �3��V>��o�G,-fyah����¥L"~�	I�:s��c"a� �6O��ܠ��>��F�TO�%�A�?���4�:�VMn���B<�J�-SjY�U-�����zs��%��?�Z�@�&�|@�E.����V+�����=:xЊFM�MniA�҇J�g����"���T�>�F?y�Ѧi@�R�F�R�����M��~����-���4	�7r@��V;T=ߨq'׽�[��r����vx�"�����7a��3;k�G��>��#����ٍ����G,����M���Q.��R^����U�fEh;�g�gA�vQ����M�&b�}憋Ġ�ENQ��+p�@d���c&�b;��f��Jގ^�WA��\���a��ǃ@��#"瀴}�%���kw/PM�j���� Ã"+#$C�Ŭi�쳣���ؤupf����$�\C�h�x������ 
�,��%R���ݡ�5vMpU�1��OK6!�f���"ׄ��$� ;����-f^*I=>֒d;���Rs&�w�~P���)ŢU��Z?jKf7{(WϪ��YB��v6;*��#l���E	�>���qw����_�U� �j�&���y�S��	����.H����t�b�lF��J-��0{W \z��ɀކ3�����1������$�T��P��g�UFTp�/v��L��2��T>��=v 3~v��S����9�spL{�)��0��?�F4�� �5㏼���<@�:5�'� ܋{����B�������^$c��)�m2K�g�4�Ш a69���ν0���F����3z����dȑ��?#�W���&�K�(>�%\߇-���1`]��nR?	۫j���zu�?��F�� �|D�o�I�*�sZ�Y�(#j��k����6z��/L��Ѻ�3�����z{�
�i�,$�A/.��=E9��V���-&v��-A�R�?�����vh��9
�d�g��;U�~��T�r,m�2���v\�BuegE�	+��3Uo�Ck�
o��}w�7��s�<X�BS	�j�wV���Xb�g�Sb�����w�r�_y�~�G�V3�6��y��r�il÷Ξځ�T��Lg[��f�fp��>g��rcM k������?�V,�+Se��{���k�Mb�e�K��pԅ����4���s���M�,D�+ ���Jm_���I`��&�.��;�:��] 6���(��	k/1�T
��8K�ow&4r�6�r����K�L�y�r���������T�L����!�(7/P�iA�n��et�I! S*���}֟qT�(��bV0d��&*a��Ρ�T���-J((e���&�mЏ�}PJ�B�򕠤�9D�s�g`L�GVmC�ZTTយ�r#!ke=e
99�Kg����DUZ��a�
Vև�������g1�P��)�w���4�0Tq/�d��S�veu���J�(���%���KN�w��|}?o�_�P&A�+p��hN(8�x�� V����@""��(ܗ����踛?��C�j�UΌ5�Io���^�g����4R5r��`D>�6ɶ��}L���Yh��I!;��?� K~�"�S"+�D����W_�HK����x����Тq#�$����g����L�[.��J��6����L'
�7**T��U�a��)�H�h���"�Ndf�ic��f>�J�wlV�:��p5|X ?ޣ6�R�7 �ͻ�cEe���\R�	\&�!�꤃N?h�%n��'c�R=��c��$���Tj���z��ȄP2B��B��pB���$���H,�8T�u��{�q3nQ�R	�EdH�a���f�HJb|�Oͭ��l��|7���I��i�*`G��)�,�"�v:���}����#�V&[z@;�Bs��L�3J|�p�szس�`	'�c������	��!u/ㇽ�#UD�mq'�'�|q%��>Ҝ���S�%R��g������Y�;Z� P_s�} �.�zȼ�I��2�֝e3�ĩȬ����y��4=�����@����6x�g�aˡ9���^��@��R�MX!<���I_2ם���%�R�wX�N��">�)g��HH�B�q�����&@:���Q������̚�ф�����:�7N����[�D���/L��W	�Z���+�p�=�$��.�i�hѰ�ǬiU�k�����$`W7� ���J@I_q�y�*�9~��=���纫�ݿ��;t�x��$�l}�_t!�:���#F��&�8����5ȤJ�+� ӈ�X��9�].��gb��
�,ݴ�����ju��n��\s�%�/����uu�}{����9�Ƨ����;|�?��@&!���%�2�٨:u@sU`Q��oA��N��
���5��.��3��y����Et�y޲��}�ҳyyg�2�G"�/�4����S�vu�y����E<�t2��5i�F7eL/�V.��Eg!�|ʕ&��A��d�`�9�=��΀B��TΟ����VH|��STӓU�9Ns��[����X���<H\�E�dDK�-�?V��-����w�S�}<���-�>�49נ��k�M��e(�h�2���n'������6�a�1V!8HJ��E�h����ۤ�B8|+'��>?��vJ�D2?ux��vm��8���γ��$��>H�H�� o�𢤜_�Q8_-Yͻc!kx9�c�a�kGϩ;��*Z�����.�rt�9ے�\�t	��,hK���>�gs��������r���[����8[.��Nw�~q� �R�e;{#���m2��׈�Mn�3T�~�R���J�R��i��3�X�3{����F�%O��݈��I�Y*��%����q�����^�*���ۗ*��t)wfU�$��14=�غd�� ��i�Ď6��P�(y)��t��/��PɈH�G��Ap��=g��3�It�&%K�Q�}�Mr�H�_#��N�(�2�ʹQ����F�˕�ъ��"�n���|;�+4�r��׍ñ�fZ����-�Vj�۟�7�Ũ�����"��(����9���jS!�OV.�2�T�|�9���y������kQY���Y�9���µ������1ܛ ��C�85��O�@����\%(�ʰ�J)�]���H���<i�yݠ3��@��읠c���e�;�T��3�p�v���:��PH�#[.��b�'��y~��燊Vc����b<�k�w����g����G�J=�h0��C�`W��Ҧ��S���j��]�x�����O�фy'/�JD����������z]`��V@Ϡ�;�-̹��~x���	�E�(�2N�䨩�jԆ�h�� �u�bz�n|�(^}hڧM�ZM������B6�c/���TP�&�|����k�s����,�(A
w#A���Σ˾�y�����0���\>�>�NY5�}xZ	 ��nT�B�!_ ��5l0k�#�����B��=�	L����M߸�R���L�Dg�ZZ|� H���~��0�/n���UCwZ��x	d�1�zs���g	W��×n���*�zü��Q�Y��A�N;�E�Q�l��#�^�3��:�"���m���۫�T�`�eP5�k���Y=yԃ�hE<�r���L�S4� �a�̠����>�����"@�_ޤ>��&pA�y��K�R�M��/&I�i��2^9#�-�3C鎤p�m�����Y7�֯���q��p�p]����(poy�L�J��s`�]�-�k��ɳ�/B��k�{B�%�'����~H$���p�C	[������pV��1�]-��V>1��n&�=c��K�d#Ts�����5������
�l9l[�B�,��~���U&�Y��/�X�����|�څ�;X���30��������ʊޣh<=�d�����Լ�-3��$�f�mA���uHc���*�h,.��-G�c]�q/j�kN�eq�X���������B�k���B��}����>�m�4!���6k�,}�a��PC��$i�M,�e�R߿Z9|��їZgޝ}FǙź�DS�K��BS����Ʒ|d*��b��=�I�NCH����_]�R	c��c�cr���ʹ�?��(�2ֆ���w$h�i������7֣=�ǪS��7iƹ�P��,�y̐���'�K̕�B�#@�Q��&���#�����UA��Ns�A�\o�{e�$Ŭ�?���\E����7p��|��R6���B]h�Ď��~ܦ=��i889>̴���t_>�ߕ�8�C����!�S�ǚ��ߑT�.�4�S�I����X�@C�iPP��W�-\=��Ԙ&���,g��_�/xKJ)��j�ҬK��~̉��=дh���7o�1�_��|�'D����M�:	�ը�	��&٩J�m5��G}��ܡT��e�GmK3t�m?��M����nz�ae�%��Pu��-�}ƻ���
�Bg��?D�����yp �/����4W�q?	��dv�h6	^5C>��
C')e2a�GeESp~b	|�[�+~7��}}ژt^�^o�������dX�ť�ϵbu��u<�Eh@� V�����P5"cU�ϵ!���lp������V|�+��X��V\���G.�`�͉j��m�Y�G3���۳,V�(�˭\���CӛW]�X~�c5�ZRC��ያ:ti⪽�P��{��E��A����T,)�I��u;9���o��$��Yڶn��r�D7T���x���c]E�6�֤�����/H^��@����zK�耔���l/�$�9N(:���P͂6�{@	�p��J���WYe{XQg))�=E��1-���K��3��JJ����uܨF֘�L������Q7cݙZ��9�m`T#S$��=1����5�s��ԍݴ�uނ FbYI�s|f�b&I�K�!�ֆ3�)o7�%Ss�P"�-z����	G���J�a��;����ي��,��׉t;G8�C�BU�x6!��P���0f#�"Wfn�-�7-�D����be�8�[�N3&�?�wR�JJ7�����]h�h�zk�3#�:¸]w׹ր�~�Q#7:�P��zOQ<`Ô�����@�y� 2� ��Pv{�Ҙ.�;��]+���L4�ls��������׏$}/�G�|X����C�+/rͬ#�vOB�X�CQ>ps;0� ��PU�܎���G�W����~��k�ʈ�$eL_��j���G���I};�5��ݢ]�(V��HcB���ä]�����,���h�ً���8�78e�M��x�ޞ&�%ZT��5�0i߻��x12�K�D�����e�!�������%� $hp,�I@�t�8�Nc�:b��{��1������h�W�||�C��T����N�aFn�U1�z�Ň�A���Ԏ���b2j�x�M�yP��¢m�U?ez�vGɈ�)��T{�l�^�R�Qeһo/Ӗ�(WV��d��iTG��@+.'�fؾ�쮝q�U{��U���҉!0�4b/KnT����l��n�_���;��K��1�DR�ĺ���Ԫ��Xp"��/��ȍ����dA��y3��TM��!b�Vs.50
��S�����
VJ����MU']^��4S=����r��9�4����^!���jŝ��oe�n�an;���}:e@OtM*�6s�Oa&1�~Ο�ǻy��=�_�Ϳ^�qupH�_w�xüXޗ����W�Y���^5ߨ��=�i�WP�n7�n[�Ш[\-1\��N���I\��BHpb�q�b"�ጹŰ�s��?=1�k�oS��^c�o�Pv�6�b�Z9H;�#�vfR(^���b�t"EMS��j衤<L.����j\P6�ȿ\�U��l��,`yJ���g����>�q�|�j�x���//�s�h��9�#O����K�]�1��_l��f���/�5��s�b1"���H�h�"�֗���Y:�� ��ה��:8/����R�5J]/��~�_��#�b��L0�:g�N0�Rj\̏,GHC�NY�y)yz0zv�f|�\����7+��W�{�4�"m##m�����*�����E�g��/���ysE��:>)D������+�P������Jߦ�y�bI�I*ݽh�������$	�V�bw�ݭM�ȷ���?a�RX֒>���WJ�|����W��%��h9��}e����cf�z��$/1��lO�TQS���yj��YM�4�OH5�����-�"�*n��|��㗃��f�U��	�s��
�[@�N�#�f��+�Q&Vd<va��O�3�n��X�ye>���e8V0���a%-��n�%aޗS~��;^k��j���)�-��~��^�}����%�(s�F�ʭɭ�.���j
k����)3Rȫ)�r����Zc�^��C���m5���<��q�g�7�
4����7lzkj>������� ώ����_[Mk��d�%����Y���F¦1��f
�����ߛ��1���K���O���2Y�<	]F� "��4��ɸ|;�?�K���eE��w'o&ڢƢo�_���iw̲���N�I���@��2�@u̧w�&��;os�q��U�Ȇ?H ��,�?T�>^ǗZ�x�4y�C�AՊ�x�]g�>>;Ǜͦ�������r	�j��U�`��:~2Ⱦ�3PXV7<�'\��j0���.�iun�<�$SN�CG�ش܆���t������Y�y�^�c�h#֦i��@�94bY*�,v�acr=���+��uAI�&h���W���󖰹`�tަ�?hR�s�jAf�Gd��(�[��雘cQχ��5�yXa쥍��¼k,��l홞����rQ��a"��+6I)�Z\�4��!�Vmo�S`+D��P�JC 	�@�(4��G��eQi�%H�Q��e'3>��P׷�J�0�,&�(6����=����b34.��&����Xe����W��\��R��俛g?�B��������� q�d~����zI���Ђ�Ɋ�����	]nd�Rb��뮦�a�EC0xUL����Z��ţ��.��'K�A/�s��D��dpᩋ6���z��[�Q�����6��V�nLR
�ím�Ee+��jl^7qcm��G�}�<�R�q�*���e��.�i�ɼ��4��I�jz����$ -6aRbł�S���i�,"F�t�/��$�=)���.�=5��BWZ�j��;��)�<�nk�.�����[��d�f`n�Y�v7:0�5�&-h�85'�X��f�x��Lw>������h��Ӛ�:��Ju
U������_N�yE��b�g�A��\T�[w��>��s�.`��u �ϋ* �S/���vYW���5*�-R�`��y�����PҴF��ն��<5��dΚ�7�._���C|��/�T#��,��9�0�熒emզ��
h�]��`&�V�J��gJ�Io�Kp�J�׹���[�#+�Ş�5X���wLMd��"�D�:�|�;�v����� s�m[G�m�1���էmU�������JK�s[d�<����f�Y��}k��~�7�r�*�ּ 列-��=��͵R�����8R�?6v[��k�����`pw��~���Z��e;Di�)�4I���0^1�*���]}�U�<&/j�Ӕ1"��@���olÆ'�xa�б9��b1�t��y|z�#�� �G�� ��GBW �ܫ�d}lQ��ll�U �Y�w�vã52` �pz�"^�\j'�_�gH��d� �0��{u���˓�����ߚ=�	��%~��F���S}������ýj�MYX�LӴߦ���}��(gl��ݗ!}1�\LK������t��&�T;�~�f���V��bm*pb �Iw͕�@jG��̹:_�2*�P�$��K~X�C�2����t+�X�kB���ۼ��S����e��9�t,o���@tlM]e/�1�f�f�s�WQ�7���/?�-Q��l�L�~k,�o`2��r0It�h,6�¶���e;� b���B�5���]��&��`�<�����$�j8
YA�\<;�!I�׹�t��A�1��y�D�he�
+��F.n�W�"�!jB	��y	__;�|7�_��]�:�H�Q0��xbn�K���r�����~�8�ʖ�˙+d�	-�T+{drkA\kK�G��͝%�6l{$٣&j���Bv�B��}��ESѸ��'VK2�����fv~z����)�+o�*�X�������rBy$�����Z���/���Y8��c�D�,t��"�-��o�>e��o�s�G�Y���Gz)#/��8���Ě܂k�9֛�1
ס���ѕB��zg�PGL#�5�A��{�u�s=C�>���}Ҫ)E�1�@�k�*�0&��	p 	mU�?��`#�%�uy�;�MHZ�+���s_����2U]Ì�H8Ճ�������H��܏���>�Y���&�c����A٣R����!*&,�����'��#���i�z��b�xq����9~��fU�����o�r��=�����|J�u�
P��*�H��?���p@�P�!�"��R�ʏ�!�s-��^v�E8n�"V�.�%�!��y2��Nl��h���( ݃`����P�Y()A䍽k���F�Vt�M���cx�aļ�n{"
�v��\~+
�BuNfC$c6�u��5'Ee��Qm�=V|b�=��GA>\{��V�ΰ	��[�v&��l:W����ԙq��i�UQ���W��F�m�3��M�(��Fc	��|�y�3U"�#�N�-���ڏ���f������ްi��Aq�����B���@=���ִ�����wuX�=�r�nl�.Et
�sE�	��[�JF�j�<QO@�c�;�(|��x�̜����@p���2����49llMG┼�XEwދ�+�\rd�J%��Y-]��L��uD_Q��v�\�Ī�m�\^�'E��z�.�B����q7��e��6!6C���I���ąO�"����9Yl9�� #���e��n��,��JN�����u����8�#MR�)�H2k�K�����bf�Pᖅ0��
�����x��8���ȉPsMQȩ�z�!�*X-�� },��E��&��A����K�)�<b�&�?�uR���s*��R3f#W���9�j�vf�6������� pf:��jDdGk@�g�Ԝ?�ϣw�qR������0���4�B�����i��J�#$pȩֳY�[�}18�2v��
��O4��#�q��5&W�ϐ���D8�~(�=cJ���T\���^HL;�ч��|ޝb�},�r+*��vm��<y��C�r�^����<"[��l��n�/��bO�J��ǲ�B&<�F�uX�O��Qwyfk4��z}��]�}_��q�y3��S��<�b P�����<�}�j��{�]s�����e���Zt���m�{i��:�!�V%���A?�3F$�<?�+S�w{c+�>X[��=�Ɂ%�չ�di/�yUgD��S���=�ƃv���wP7��w�fj��e&ϙ���Y��z4���@}Ժ��E�~�B�b�U�6��&��\�����b���E�c��Ї"�	��(����& j�!JFo��h�-�m�MB��;8�{Wm7Q���\��N��6
���s���!YK�@߲Hɦ�߽*����0)��D��G@�P�i*�k���<%�5wYIb{a�z�J=d�U�l�p|xN���g}F�¾M���}���_��)��d�9eRz!W�5iAΜ@��&�����xk*\
�u���af�KK�W�S�S��gT۝\Ok6L����z���3M-�/�fN4��5xY�񓿾��7d>���j~�Y�x�$t�=^��ܯ�M�r_fT�ov[@ܢ��;`!�����0�?�cm�j�kGQ�o�j��$�Q�X<�����NT���o�D�e�H_ɟ`*7�^���Ic"\�"�=׻��6B1셔�@0%4zgJ799����`����C�= ���?=+�LE�\�k�ѮIҠ� [=�{�����rȋo^e�`Ł�����F���(��M���~��m�q�Nȵ�-&a�B�O�_��� ����)z�٠�P	���$�?�#tb�G��C�v_��^�͉i\�}�AS�)%k�G������E�۠o�]ս�&�:x���$��gXÿ�hY͈�@j��[�<���50��DܴCc爈�L/\�
7�� a?TVrd�I�R^�x'KT ?80:��BP�cux����ʚ���RD�Ͳ���'�7����)-`�/�f.���ðǁ�ph"Ҽ
�8ur��m��[~!$[�l�Ы_����u-}N8�8�Iw���vSCq��g���X�������#��˃��oN������B��t%L���������Fu�K�=��σ�*O�m�/��!�꼈�gD�U�Y����a�۞��;�U�:����}����qbZ���=U�U\�Ż��k ����6�Ժb>��x=w�C�Ƒʲ�z�?%�_���d�T����*�߿,�f5Vbe��{�������Uw�v��UQP��25�mr��b��Fȵ��Q��)��[�s���w8*�[1��[q�-���4#HݠԐ��5A�,,�i��)�@���FD�[���.���s�n�o�����Z��R�F��&�a��v��A_ �K�~rFL�7�����kb�7��P��0l�6�������魉���m����Gd;C�!cvlbeM��F~��L�QvD��A��d!|F�y*�0IOA@�=��;�Ϙ�s��f0,��d>A��s �� *��C,�K.��%������(k3$WkO��پ��� ��;	�^Ӻ8&!��������a��5I����g�36-�;$��{��$�`v��P-ı�/�ۏc �g�q��9���Q�V�o���1��.��o9�3c�.�&�go�,��5�X�0`�x�j�|�� ����C�U�q�N�_m&��	��ř�"��ʯu�0`�L@؏�R2��:����B���D�I;��[��B�����')�:�y|��X�/��6��H-�g���ǱS�ɜ��^1�q-���(���f���ݨ������t`�+�_'���U~'N�K�֭a���鮈׬�(�=6����Ma��@5w���#��]�}������sD�J,e�(Z��7�Вށ0ŝ��0���j�����a��?��2F�Uc�7�v1�5�97�~ܭr��2�ִk��/P"��ͫ��]���tU��ىڻ����Rc���>VvL6/T8�A����x�����"r��a��,��IDńac�8��M�=�D@�Z�y�#��Q�ɠdd~���Ɠ)JkQ�C���s,Q�����X��^� T�_h�����Wsڂ��0��Ԋ�����(�B��$~>P�F�m,���0�$���s t�=�[�м���%�L�^���������H�ɱ�B�)�:�Wm���Ѐ�s������� _�}s�Xg�'a="�o�_����L��9`X���-l����po5j}n�izi��_c�@���Ҧ�l���F���?o�Րƃ6
��8���[qӍ���O)'���)���x�ݬo"�~'��:�ʯ���|s7��7�?]��ȱ��|+�Ny����׳ϑ����O���9�j�O�M��Bd�V�G[/��j,Ya$��	�e��	�����G4 ��]�P�I��g���f��c�qQ+oxR;y�ݘ��G�-�͛��o8�Gk��6�<�2�X���3êBF�����vGdd�	I�X#YZ�A�y{W��Q�v9��xHM�)ӵ����"y�����6�z�G�,X�<l��a{Q,a������գ�}u���}��B�֭I��/Ҳ�)u�#p�M[S�L'iB��OJ`�M��F:���Ũ���B����~���� ���$�Fn�u���31��?�&~�,)Y�j���>��/z��WT��-���K'Z�3pFT����܏�H9w4�]jm��1͝tT��������犃�����j`�8�q��S�]^}ڕ3Kx,A#կ$�c�gyu��]����r���(f#��KD�q��',>����$���+l��){&�[�;f.�(5����nȲ\ן`ca�ѿ���k?�^�;�q,���9��ʐ��q�q(�P�s��\*~OG��,S_�=��}��-�j�`��T�A
�'f�G9���g���cL�@,�sy�(O=�-��:���*��A��\��U�]�������?�o������ei����f���Ӂr�bh>�}K����{�I��]&��l�=���E���`�_�{S�g�t����^2��m�Ͳ��!f��� ��H!AQ�2k.��~�\ �x�2F��FX�[k)���}�M�I��G�u�	�-��!ke��)6 ]�� �/���u3�CS�ɨb8�N� �R�����\��5���|�橌�c���-�U��y�����ˉ� ;�8�+X����d���v�G��_XGøM F�2+�v@��Ә��.]�eCﱆ|j��3B��9(�\�n�����	2ų�c�������zG_? h�%�BkB��}����v<z�r����c�ʀ^���G[o���wI��Q�W�1u�
 c��n6>�G��0̩5p�X68��)�Q�`���-�Rf��^,�����SC.�����J�⣯�mɇ(j�`ѷ<�t��ɼM��m�~�LE���Z�f+!+n�pC�>jvG��k����G�y�Z.̋��I�����KK��-j�
�s��=��i�ک4q��� �����Գ*���=Us>㋊����/H~�/�/�k�ϭ!%��J��yNf��g��fѫq�ζi\�v�^ (���D��N7܆���>�����2��qPHX٤�ٳ��;�`�":��'�����xM��1�O�h���~+v>��7$J�j(U��ꄟ�}����V7��6��H�1����8<��Y��H���Y0�x
R�}4�h�s���5�V�3�&6"ʌI��>��y-����2��1����*^h�J"y`�rS���?Ȓ7Nk*^5���jAl�:s�_�}gOH5��6��F��#� �E��%	ގ����݇�=����p��� c�G[�޾�Eѐ5�6��_)��G=V
��{P����v�)g�5o�!�$ϐ1�o�R��I�~U�T"W���"���DƂR�
Z�[�w��w_����V�M=D�(XpqJ�"T�*m�gZE-�c�a_2����G�Z����*�,�P���}[�:��*�?�����tŅ�0:�ޥ(�v<���O��r���*��̦]r�E��{XOej7y�/��eH�XZ�\ڂ����`ޒ�>H��p8�E�O���+'P
���Ώ�D��Ž�O�4}6�H�+��o��r������=js��-.74IT,����Yy&�o�c�8&#G������
���r#W01�=�[����iʂ��ګ\3K=5��ɮ���O R�\@�o�4���B��J����_�c�I���:�X�*�F9kV�i
z<i~Zr�,b�U����)�SˎNys��(3;�*�GH.�����i�vp����9|j�#���)�B����4��)�nR#���W$_N~=�u�(���K��;����Bs �k��J�"�2-�m���A��{R�Pkɨ��	R�0���k�J�qό �Vlo�ý��>:��_IϙS�8�X�:`����gz������ତ��TD����)w
 �%2�ነ��
���	'I�j����-;��t!����	��Xc�F��� �J؄6���@�7J-<�H6�Z��b|<Yq�{Qq-/�7t�o%t���Mz�J<��$P�l!(m+=gA��ɮØ��ҵu��pҚˀ 	�͇m�/u<?����-����`C)�t5�uv�^|����V�`;v_����b�-�d����i7�M��\Wo���v�V`�t�G�_�O���H�D�a7R1j\�.g9[�??�{�I��ۉg[�gM,��=�|��z>��������(�;U��Ff��d�.�_�r�A#�,���;5n@�N��n<i���\e�wk��F'�w�S��IUt"/C�~V���
�НU������>����r:/,^gPD���K������3�E���j����]��Mx�kq���r��O���X��ʬ����6���L�q0���E��1������=�Ъ4�
8D�T9��Y��)o�z�y��<Mba���O#{W}�V5���j�?u��^P|�]�^��U	��7� ;lo�\7�ԍV7��H7�_�K�OV��c/q{|@a�b�= "9	�w[,������Qv�=���C��yA!KSK���ڭ s�-���2�y�u�wV��G�ך�j��9���l��l�[��	������:�/R�T�/vj�rp��آ��I�$�1���2�<!������ۉS�|�jZu��$!O��J9��MN�;@䒹��\?W����E*"WJ�2��>���:�y��/����ab@��-Z��+��v����w�h�wLS��]� 3WTV��.;�Q�$.�pk�������ML#{�����`��b,R�@B5������_����R�o�/���X�
c@_���h��OP���<�jq�X|a����AK�I��������4�>���n�]���� ��]�%���Ë>�0=�](V�4�	+����5��Ӷ�x"s���kTp�;��b��]Oe�1ņ�MMn՜i1W�-��1�B��Vv���(ɲ��-�W ��تN!Oi_��r/�� �D��H��<2���(�g�������H^:1I�R�e��B��|՛����jL�)�[�8�d�kd_~.Ɉ�;J�PJn�Y!3_ݜ$�gX�[:|X=���Y~|�NȅN��EM
(��\�y9��D�����_B�B�e��X��$�ACP/�(O�mi�̗��g��Y�{�(	�!�I?���Cz�P1�j��?�̭��]��s~����d7���0p��?q]"�����{���6TD1.�@P���C���37N�8|z�qA�g�:h���l	�C�]s��k��/�+3�D^0W��K����h!�M�Q��U����$�>�!�VS�z��;�_n�~�kf[`d+�[4>�"Q�2�3�c�G���1^�^`�k'<��ȏ���X���,����"�'{�!D��r�Ϫ���x� ��֖ݥWt�m�ߣ��5���bY�E �kLbÖ1+�'=��P^6.�o�S.ϥȥ����9E�}�6:�Y<��D� �!�~��'.�I6&���C͡6�B*f����ɩ��g��:i���c�D�q�_�&��j��n�g���G���l����5,?����tԠ�4ڒ��:�С+��bG�� �"3���g��9��1T��!/,֐��)��,tl*��Ʀ��p�U��{��Hs�d 1VV�~��Z��]LKX'� �V_��W��u�~��2z��<9�߇���N�K���DM�Q�q`�,��Ey�om�k��5�����z7��B�s��Q��̲zJVf2��G2L�pL�"� ���`���Ȟ�:'��vS#a�8-�a씞����.?��N��Rf������GTA�:��.u_��������[,�~�j0$T~ht��4���g�7��E��N�+R	���̗�]��@.��(�޲u hhYO��g�N }���F7��w�#�3���^~�>�\�8�|���I��K�M^zOs�W�d����,�I��d�vUT%��9���0��e�H��v3���%!ϩ�8|0Z7����-��7�r��l�,eFԇ"_
��n�D�A���sX���6�)�qע�&.������ڰ����Jb����\�e� K\T��1��%A?s�����zqXx2;�U���.�>.�������������a�m�N�u�J��4�.d9�M5�ʉ��Kr�p�*����&Y�}!K�� �]^�Ä�Ȫo�`b�M��T[)�GzV�D꣱n�I�R����/�������
ǉJ	"vI�]᧶g��j�۵z�b����r��o��[5��tO������Y9T�S �i�G���i�ՅPe���WoGw�ho�i{"*��o�KZo��8�L؜�Tn���Լ�YSh����S}���sl8��n��g��cPz[3\&��U�Ux�W���4E��9��AqlX��xD����=#�r�4�?ϛ����p�X�F=�Lkٿ���F��v�AFO���G�u��Ke�7���JTA|��;G�čv�$N˂>r19�Mq���!�S�F3�V{Z��d��I������+5W��d����9)��Y���bE8F����JU�2-��@U�3��j�����F&�Vr��J�ZLX��8�{nHCV^C�j7�W��(H���j�ԉ�=��4F]���
(��G�y�~	�r����8���e���auc��Ӷ��H�PȌ't
�1Ɩua��@}����*KRj
��%�/m�e#�Q:7R�a4�J���̻]&�6�2�	�JI�؃�l�FH�ۛn��r";^~V�Ρ��Koz��7
	���w�)��W��tR4nP퀶�G8����9R�J�m���J,Mw�7!��K �h�s�����r��Wʈ��rf5槲;���8��_�k��;%J��q�'�o7g�J܋��s*���x�iF/��C�vEA�z��;(u���~N(
��B��!�ې��s)��(�{���%�2N���������D��K>�3ݦ��JԸ�U�6����/�B��x;��:�;��B�G?9Bzx[�-՚t�cT�p��Z_�4��"�V��$0續d��Xh m�|�<�r���_�īɺi�PM�0��00�#�2��j�|�@��Q&��� �[��r�Gh�gY�~e8�o�^��g�[�Y��<���r&���.�r1�w���W�+c���,�F���!��\h)����Ӧ�_���o�J���DgW��/���<z5�%�9jU��� �ܤ-Zj�8[^� �]
�R,��O/\0�c�@���k�����˞�Oy�}�?F!��5��Nٝ�j���6�*|���D���@��(z !��R�bW嵄CR;���[������ɦ��~t�t����8�+$����&��jp����+g�tI��{�қG�O����5_NA��|���`�^Z1��{���p��A1x�,�n/�k�9�{ub$�Ya��6�9�a���"�]xT�c�Vp؍�uSm|�D�[\�V-�.�0]���tɺo�OI:����{�t�ѵ�L�e3��E=j�d�#Ҁd.�`��Yk	��m�z�#���~>IPʌ�Ö9H����a���I�HZ�D�%��38���Ei�R��[c'Ĉ��	e��!n��M�6���2X��Y�O��hH�웁�*��M��8�a��W�����x�%���-�r�O�5a����6~o�D2�\��N��%�	�OI�|�ػNČ���f8\!�G�R�+�^""LB�Qy���^����l_���(&^*���Z���LMˊ�Xr�!a:9EJ��#Bw�bI�A����
�+�(s��c+5���C� P���%#I���.�p`�����m�$�*�@�T���ⰿ0}!��&��I��nr���'90���2D�,`i�\L.�IjX{*	���s!�%�pPsH���Q#;��]߮�[I�*��v��Ba�(L��~�S�~�P/8�� �	�j%'b�J�_Z�d]kb�kY��o����2$�=j���:��,����v �F�����T2����r�($w��e�I�`���u[]T��7g��g���� 6+�蚪��X�:�q\�#�*�t�R�(JN�q�N��+��*�X24�뷐U�M��GJs�2�ֲ�����b��eS\*��P�6�)�k,��x�=���ў+��6�ڗ��l[��cx���{�TπQo���U�p�Uж[2�vDl{��MX��q��uC���|�7���>�q�\m��\E��c6���go��+cg|qETY�	E�.��V�f��x}bA�ki�]�b@�q�w�q�i�6Շ�Ո,Wv����N>�XQЪy�@.|�K�*7�+ "��m/��"��y(��o��H��]��Mc-�O���7{�9�Sq�����D����},��Y2O9�$3�m	����_V�ɵ���D7tE��1�;��#�E���Č=��a%t��C'!T� �0�:q���2*e�hOG��8@n3J���mI>ǥ���v)���0�@�����f.6�>'(]ۮ�d��#o/"+rUd"����/���N{�.�E&��X:-6��]�r��_Rr��$#�4��e�@ViԴ�%P�"_���)v�E���6~�)�`���˙䆪Zͥ�B3�h���:^}��Ndʱ@��`~�� k�M��s�D�������3K���vL�� + �F� ���8��d�8)�sui��U���;[����wX�ވ������T�ge�E֖�s�s�t�1A���4w���S*��<-q�ãJ�Q��Ɓ[ˍw�8��T��g����o�7�T����?���W�,���]�o��BE�dHB�Nt�G݂Ξ����	"�
���3\���/�ڠ�Ɩ�a<f��|��ڈhs.q2��SwL7���N��0YmQ�]���h"�; Q�3�����jF�M2��Vk˒�|��>�j1����B�`w���[��*�����=��lm�l(����!� XL<	\M2F�}p��qG�ۢ5��Ǩ�����B|�N6�
�6�|1d�$s���c�l���@D>`d|"���H{���\x0��V0��΄d�䎛�h[���	G�Ɇ��[�eiM������D�x��9�9TTD����:���j�A�G���ٓm��c�S���0~�{͆�=���P�,�R�$
�p?�������]���]�B�њ�*z9J���@���d���S\���b��F�z'2���ǍЫI5a=�u����C$�w"���l�i�ww���T�*���Uo>`������cv��]�|���J�>�kH�_�_�����1ו��P�
��&ƯVmB��te�<�6%���#�G_ ���nc��hz7�t��UeǮ�g@fn�G�pL��.&�XFu�r+�Ω! 7v�<��_�2��)��d7�z�cHs��(9g����t�ظ|C%!NJR���c bi��s�^6ח0�HN@�����C
% �eJ-.2���P�vǯ���G6��$���]��ܤڝg͵L��*�w �s/�H������5ym0#ޙ4<���
4��P]����U��[�5M1j�7.����5F����%��9Y��'�|{���%���Q�\x�w��|�b�����r�=�X\�q��/�;�&3�ㅇ �T~z��0��[�ֵ��iaI9��O!$��GgG�:�,�M��<�bw��䰚O�ے�%��B0}�Β�o��Ӛ�z�+/\�����Y|�5Q5+��I�Ǡ�Oy<ª���ɢ^�k�ĭ�����ȭԡ�(�<�B�&Ė����=��I��ehJ�cy:]J�8��<�/4,e��8z�Z�vMR[��Nb��.�p�� ��0���%E_k
/��}vjn�5Rr.%���"T�]]�d>w
��7��i�Y�F�Z��c ��U[�j�~a4#���H�ଟ9RvM��5��N�R�}e���!���k'pt�Ds�VѺ�%�N O9�A��Ԑ3C�������ad�T��T��1c;U��'�j�:7QE0ݛ��%�	��kh� t1��16��ƹ�bw�>��_�w{VRKD��\�,4�3���|F�J�,ע���:~���qS��˾Y1):�
4��F����9v���L��qީ���0۫n�榻�}v���u�[a��1��qϢbQ#��V�-*:!! �������V���]���ydl��f8m$&p/KZ���x�(dqA_�~�W$�IIVt���N���Q�5#h1Dcky��gw�X��8f-���e�R�6��ڸ��)+R�H����vܡ�A�:z�$��[]U�l����K��^|Rp�"���=��h�e/� ��:���.�����$3���}(���������9�>wſ	��w��?�0~��w>\��"�y �v�����6��s���Û���hj����{פP���N���'P��+~vj4�Y����>��P��g�d��c۳��9�t�4�gu"2�+r���H>B�yr^P�'5��F�w���C�\�	C�=)GR�X�tx�����I���й*�D�O��A�:��;�W���� >�dNNuH���4�hy;�w�\RՒ�@�9��������uV{���~[�kֈr5��,�VjEO��\H,��R��_9���VC6�
c�.��r<���m���ar.�nƲ�	x�!�qL/J��X�rw�v��#+�~+w���uo�E-�� y�#^CY�r��7���qo|��ղ��aC$�v������$��]�+���$�.�2��*0����Y?�"�Js[Ϩ�Ys����αk��1��#:O�9r3�fzk]O�_�H�j�3w,�����EݹÏ���/+gS�� �d���3{�ǋX@�ν��%� ����}������䶉�,&�W�DM�Y�$��u2g�3�p���.�>���,��[�Sv��EU�i�RwmGWX,Xw����>��;��yV��7��ܸ9�NB���E�l�OB����������q���: &����7�듣ȴW�d�$¤�m4f��	4`�ސ�\�����9��2���!���OAP,�o�^��*� 2o��i5����K��ߺRnר	Y�T
�h���ճ�nD��g��)�V��������@7�����-�\Ō�W����+%�K&y�*�dw/wf·�ۼ��=��P�ݷ >�oOu%�:e_�r���܈E	eb4��P�C�� v�@�� ī\E����
��V��&o��#gz��O�L���wB�˄��vMG�*O�o��	����&��Z�3aǃ2n �ȤYe<�mX�S��)�z�[F3������%k��g��c���f8�P�+�v�zh�E#1 C�g�s��(���Y��L��L���[5�_8�!_���L��/�������<�]�sj
��΃���qw{�1X**�y�6&��*�������	�#���/uV1�>�yW�5*0��ID${��41W{O�SF�����cĕ��R�]�x��{<�(�͕z:Db21�شlӛ���"�e�"&Fճ�g��`�#=�����|�_�F�DrVT��۫�oP��Z�g�][᫄�w��xܳ��<���#&�qB�9˲���%�X� �]�Ήb`
WkO'~N^����5l�GA�V��d��
��
v�qZ��f���%�\�/���0�搌~N�́Vkf����F�A�ߖ$5
�^~H��8]����B�U�/�����c�n�F���<���	n��v�-����&� ���#Q�NG�$ ���[����[^#2�w���i ��PG�R
q���V�"&m��Ӛc�e�B���s�P���Wɉ�G M���W,�4�� �J�	%�*�7Һ)�`���#�%����)��� j��1�1h�_ʫ{��S�M8�46�:2����_[�I���d��,�1�n�s�C����V��'/�a�,d�����wD�_��{ٰ�3���!��n�L�V$q�� �:���D}��HS����{/q�W&���J�k/��JA�i����00��c��U7�������iF��Wh�x��j�#Θ�q�[�Tv��Uݬ�W����x�$�څ�b=�ʹ�����ߥn�ve�;��%�����5t�1������f~����k@��k�J.���j3}kA�G�Ȉ֌ɐE�s7=�o�0]*tGP�MM���-yכ�T=d�����z�W?�9�������o��wa{��%�耡�C�r�G�Ws��?�Z���^�)_�HvZM�F�U�d���0�۱-8!�UT`X�S4��E�"�Y1�������f����eFC��Ohh�d�h�ּ�� �tj*�i��/!����-*DC,�@����(��G �2�V!��<��(�G�N�Fn���ro}@\�Z-W=��j��|c��{��h[;u����?�50�#�^��v����*�_��Ѿ�&#�t��l* ���?�+ԂOt��pӥ�I���
��Z�������e�I>1�����ԉ�a���u3ǈ���J1Ì�6U����-���P"�%�	{�G�t�2���Yã�JS'�o����ބ_���c�̈́�d�<+�����t��b��Č�Mӊ�2�\��N���n�f�!q��M��h�8���'��Ϻ�D'��d\=G�]�L��{#=���k�Zh(��5Z/���m(.ͥT�ZR����*2�=��8�� 
�&��CE�~�'r���Nm[4�[�����iQ���d��%�zI�H�^�����_m���B�X{�'a�T�chf���AЃR���K��/�����\U��Җ������:K/���e�#��T�wܸ��J)e�b٩�����r�J�Iϸ&*;`ЕM{n��L�qX���8�q�$A6I:X��'2sX�p$��Gm^� ��?R������p7&Y���kjB�\
�9>f��~X���`Rv�����dp߯-����䬄gͥ\��
ӥ}?�FWR�w���������~#��h�*��h�m������2$0���:�<���V��y�5��O�Y�.�&�Y���H��x��J�)XTᑌ�I}_&<�!�`�H>\��O��t>���<�r��;����T�1&�+�@_z;[��\�H��H�����P秿�j����dg����0�߉��� �<I�)p{9��T��R���u��ɶ�[�J�*�Q�D"_U�:s����.��9#�S)��hDN�*=2n�g���t� p皲�����Ľ�_VW�#ԝ��;el�%�E �������t�]��Bv��/o�~[�Y8Z"]	`�G�R�������@�iWKQ�Ie�KފL��d��-|�:+�=��U�tKm�T5W�=�y5ݢx��YР���
5v�t�QG\��]�� ���)V�[��V������/��"}�O�/��<=�d�@��!	���e�]B� �8��a&�m�ȧ,`S&��ME��x&��Ծ�V.6w.��]���R��03h��G��a�sNԹ�9�	�20
*����'���{�uD�~vgYq�!r�g�_��BM��8�1U ���1l#��0K�&}T�zp;��6�^��FX4�-i�>��p/y���,�?i\w���1|��Npw۹U'����	�u�y�FT�'�6���(1�τ/�7���S�)�=��^�8ټ���%�ӗ3)E��E5y�.&��������o �%xV���|���u�z��5)Zc9�j�kw����ĽB�F|��5�vId��JU�����M��!���c,MX`#.�H��s���������]�� EH��y���HY�����q���\N��|f�A����'+v$�L��������P���)F����s�����^K��XVFR����O�V�լV�o����#0|��S��g���{v��֣��k��w���L�b��A����_�d����<@�0'7Q�H-YAkf>V�v�ͥb^E;��:
H]���P�ъe\��H�{�]�t[�5�o���`�ǖ����Hr���t�C�Ys]��N0R�µ���v?�Ɛ5ɲU������A�2�	���7c�*��^LEo �a$����i�͍O���C�V�#���M�ޥ��1!��k�Z��O�6�,�@�e����y[�2̴�L*a�fŭ��������_��ӣ��ɣ���wŚ�Ϳ.1���Mm~w~kTSc����^K*R�V��z����eN��r;����S��2��mt�>@��w%��9��;#�g=����.Za������\T�����jp�����pʦ�l}�����J�L2@+����@�U�.{gD:}:�n9�g	r>O������
����3A��Iѵo,��l�5�ה���ɳ�>"��}q�(e����v[wj�P�������h~�3���'�d
���K/�;o����i��y�����D�P`�����m�(��j%JS�s�hU׬��� Zu1^���K��L7ZFF�i�C�7����y/�aӿ'Մ�N�=?Y؉v�f�0����V����q\�H4�I!� $�|�<ہ����L��#bI�V���ٹ(��N/���l�I%�?�?����5�ǫ)D���7�#�֜��Ϧ�d�����y�������_݇Č�����*�ٱHIJ�u���1���Y {6˒�&i�/�~�-�<R&�����-�ʈ;���;�{$y�9��WR7��o��X��yW"�4���VN��2��)ګ��I��G��M�l'I�H޽�Q���r�T1Q;��\�&�c-�]�QU�I
�>��r� �MCz��LGR��b7�V��{7=t"�޽�n�uг�=׌nq�5n6Sk%�ZZ�7qY��mN/D���P9
�{۰6ב͘��F��n|�P?��i���5���A碲�][�²쁴�s;YPއ'�&qh���j���Ƌ�f�I�c&�ȧ��lL�Q ���w�|'n}�#t�ȏ�n�E,MOp��̠�7�L��%%�=NŰ�ԋ��P+�~�����}L���0+ݴ���֒��+���1N��/�ó�ݼ)�c�.�FY��i(�)ן6a���l�Bp�"1�]A@������O$��s_K��0��t��.��v���- C@�Pm��=���d�-F�.w(�~�I2��7ȕ�/�.���N�p�^�k(Q0���}�׊FC�˾IV' 4l��;?����Am@�ݑi#���vRK0Y|]Pz��`�#���1s���Q�d4!��{�8�[O/�ߛ
G�L�I5*�H�V�}�1����e�N�e����My$5��#���M��p?�QE��g`/�5��'�n�oѣ%whj(��{Uq�#�3���g���v�Gj�r��}���_b�Pl��Q�͉&�3�����6�OzB�i�鈳�:Ю�F�쒠������_��.~T/J"��SV> ��Pɂ���Ӓ�A�Ů+�=�#+gI�˚��&5'}�������'|TUm���L�K�
���GcQ��2*�'HS�QR7���4�IdС���%'��_����'�0��n��Cfꂊ?&�ˍ������g^����!�>4AU��������܂V*_�C �cͅAw��-&�)#tR��8�[o!"����
�lÊb��'�R�jϧ���e����w����m0>r\�u�[�{V�)7Õ�S���WJ�g-n?8N8��I�&�i��+�c��Y`n��r�*GI�J���D鬐m">{�S@:Aq���oQ8���
�z�^��[�Ž%��h�[>#-�o��@��B;����'aD�Z����@bp��tT�,(����L�5���__�[�_F�𷋻o�J0��1�)m���X���Lx&M�b��ۜ$����,�Z�[[��=�:=��ٶ����b�i(�(y�=�VI����u��oXS�>�t�֘�&�?�+���i�X��*��t�gy���+�E��I�i��.X
��1��mMG��X���MIHd,a�;8��s-�����2�
�l����`�_��c�U��@��C
=i92��3:d�Qc�b�|pb�)V�����b�Ɨո�kS(�s��^�`z�Lme��|1�W<c�{xu��:t�e�H*�����N�Z�~
	���4F\���Y���q��!ϰ��0jF�І�s�Y$����i�<��^��i�֯����r?�"���݊l )h৽�R���(С�)����5S��&(l�,/���푩[dR5�s�N֏@��Cv8/����\�Q!�+АP�H#�l�d(�)����&H2�_W�7��J�����zt��}�5W�j���b|&���ܱ=CF%v-����\<#� ,�_6��jix�E�չ�Y��#�%F�p&L:�K�T{��WP�=L�3�𢗋{�g��t�[C꟰��v�|��r&/,]HY1�A���?I�L��~�e��h@�k���1�$#�~wL�|��w
 ��-�w��6 Io9Y�(��8���eU�ԅ�K��)Z�+_���+*��y�I"g�1�9\F���v�a=����Jϐ
UX���,�z	�ȑ�P�d�\a�~��W���B�')E!-:�;�A��79��y�V,[O��r!?م���04������c��Ԭ�YJ��Z}�|��D6���қKP�8V�08I�ȴ�t~㠢o��F�Gr0c �7$�U�}2h�}1���9�5Q�mb�,B�Ӓ��ך���Ņ&����{& 2g5{8[��fZiOEG]�pӲv�Ƕ��O��yt�ď$��������+bw >T�x�x,��s�J�{���ao���!X��3E@�Ь8�Rd0U'�q2��Hc+o��;C��a�I=�t�q��:��[��2ӫG~y>v�`o���4���*�6\OUHf��r��i<'	o+�]}�t\�((1=5K<���Y��;��vW�lM1n�t��f	A��+��F�g�+@B0C�I�U��38�s�T=�կ��)n�l�-U�x�UÅ;U�ң,#�~��aKLYt*��O!%�s_�d��w�2�v�jS�q����ɋ.
�<o:���ϲ�/]��Y��Bٽ�ׂ�{ �
N*�E�*�&��H�f��V�0 ,�R�b��R4��O�:�}�C	}Q��NO��$���r��f���V`I���-Xi+��zA*@������@#?�rGE�{E5G ƮvPY) \+��h��<�����ZIh3آI�O�c�I�VH����es�"�3�����^۩B��w�	��i[�J��66���y����OȀ8�yBp"e�\�����Ц�D�7w�_�}����Ht&k;X��T����a�87U}����F �2�A�e���?)��{|�38$���~m�M_pS	Ҿ3i�c0�[��[�e���n���]��q�f�땴�S�x�$�{�-�Q�<����.��}f�dvw��k����1~U�!��}��
H��-�J�"
}&�W�V�B3�XNd���^�yp ��Z�*��W�����Y��(�U� *��XՓ#�����8�u\FEV���SH&Wk��ۀ_��:V�a���R"2��tS�a�b�8�v0:X /���˅��d�A��-����˛7�w�/�^�p�M�׃>���qlw8�Щ?�#�[w���i֮�?޻��Bl�C�6~��~�6l�0���l�W�?XM-���,�چ���	OR ��eD��sUb9�I��1
(#��R�F��_Zጨ�P�-X.�ҿ&W��.x���G�ĕ曤�q~�|2GJ�l����������"K���FE�.X�x�:�!�aX�ǯ�J\�%c���vJ�tgth�`�i5��vUR��i�Gh���Z��ur/�a���5��x�h��؍�mD��X��̡�+�ۊ|�j덦Mm���H?%�����S���H�_zX[u'�M<�P�>׀��ja�-h���Z��S��2S���`�Z��h��AΫ��B:�-�x�(\��ɗ:�����ϓTI�2>,��Q�/O�/"o�����+^��,/��e� 7�����@M�j�O��6�=63pm���V8�[�b��y����c<��'	?9#z�;�{Z������
��DmO�ܒb�?u6�rC]磔n���Xm�sଙ�g������R))r[���#�z���ۈ�n��e>��"Ŝy?������DN |�Ӕ7�9����[�SV��G�M�U{,tK�1VmE���xF+�%p���`�s���y�!�E5�R�'Ǖ�cV�	�8�tb�{�>�>x���:���tE�8�I�by�}&%����6K�@�f��ZRǄ��k��"$�BxIG)��4ﵵ5�a��^!�q�TڄTْ�b��eH��Q~'��f_�i��e��=٘O�ʠ��ϋ��t�'_}n�7/-�#��ŷ	r�0K���c���w]��ج�6Hu�d�������/��&�X�ʍ#�
w5�!�RV{�_Ej��P)-7��ܹ�Φケ�P�)i_A�@�gm�Wf�8�n�' AڸT� �([m�I_Q!�"��⎟9k�(��ɛ���[lM�U%��q�Ta!��McẴyK�`u+&���h.�a|�&sLƶ�ؔ\���J1��?���q���j�����͵�r>:�)P��)�Y�CbY��̋�]�_D I��c.�&����."�T��|���C+A�i�`'s�~7w��b"y���t0�//�!	����-kı.b���NL�֓�� _���O
��SB��}M�K�?;J�&���:�E��p�X O��+�U��{ẻ���?N�`�7S���"a�j�AƮBc��w!����7�w�O��
11A��$����
f����:Ȋ�G�k����7�������^)-��<
O#fm�����Y�u��-	��_���������S����g\@:�C�2 ���y/��]\,4U�z���W��l.��e�ѰmcMRY���_f^��;C�=R��e:8X��tj�����F_�|ҘX	��m٬��[;�c��y������rĒ˭"��Є�̌6�h����,k�w��W�A�G�{������#[����P�6ޯ�4i'D�{f�*ڵG�,pՊ�ʷ0�c?�&�RXA�ySm����9�)Z�1q��-l<�H��D\�f��\��9��Cr���iV�!j���Z����P��,z@���\�������(��"��HU����k:�����RRԹ�ų��uZi+��Q(E�`�+U���o���%�צڨްկ ?c��p�pϷ*g�
� 3@�i��	R=k~��X'��40L�����H|�<in\>̂I��Rv���M��-�j�@� �б���H6->yU�T���{XH%���>H�\��J��N���+�|��B�2̈��]`�Jݘ���eP	ɷGՔ�4��w��t��v��~B���nI9���>��՝�S~��uM��v��:��C�_��$�Y;��HF�׌��\�LԶY�������Ps�ny!����I��h�p>��]"P��SA~τ��#���L4�bPq��O��~L�3Z�5o�����K�J�Ju���_���(�����;��ar|D4��iX
���.[o�o?yj�^(1؀7G������+����-�i 8,pG�M=�t��y0�	гd�-쭗2�%��xgO��P��L��.��qB�'}Y79����V@����<W���ö����yNo�d��T��#ðF�v����9�|>
W��[;����b��	◛ ����� aO�z���������tD��a�a���P+�8Wo帾�G�~����_}&�w�Nz��ʂ�!�7��Z��"��:����	%�U�L���l�+c[ �+���9\�[
6��G<��g8����u׋Kj�1�Ԝ �����4Ր��D��35�������n���W;PU�q#�|O.�Nt��4�1yF�l�ĭ���4��8ʤ�n�A�Oң��ܓ���dC�L����8wM
K��o���	��A
�)]���ՠ�bm��W�3�u�L�S@�\��gU�/	<�����_X�d'����"?�{0E�0��+����L�K�F�rX��U���e�Gh�n���|S��O|$ܴ���A�� $`�H2��B����E�Ά)=�ީL+1������k;6�6Z�r�p�W��*O����*�6��2��ۄE�-�4��?������D;� "bY!�[.[��Q��UU�w�.`��Alt����7._ܤOMp�7�Q��c��#�L��䠊�Q|Z �����������T���Ϭ���U"�j�EP�����	�0?�ꢩ7o����̪C">Xp���)[@�r9��p*4�R�S>��5as�B�QP���Ҧ�}}��r Ss��gu��N2�#��f���|�^2�j�iV���mf�U-��I��R��hl4$*n4�Ջ��S}��:�J>IhӀ�Я!�Î)^nm��|�GP}��!A�"�� ��>!^��@�q&wMV������܄��*��U�i�T�[��Q��ם�y���Ƌ��Hcng	*eø^d.g���XW^,�.I/[-���\0�ǚ��<!��9.o��دrB�
���i~���4�֔s >����va�;h�������K�޿Dw+��i����C���a�<���Pv�����b�����N��gD����7fē�!Rϒ?b��R�ZzD�<���_X�V��$zK����X����J���O�߄�K�"Eb����r�h44~�,�f�!w#�����zi,)`���;����tB��Vg��,���,w�rs���1�wn�M��o�G!h؛�B�	��q�gx��۴����sY�v썋�kk�}��tM<�<��^ʢ�qO��{!�o�X�������]258�l�d�����&ep���A��ܡ�=�t?�@)��3z�TWq�@�U�EX5D9ADU{�:}�,ǥ:�`�bGXQ�Ғ���	�����^E�!��
���x�0Σkj� IٮTiC+}�A��Ì�掣���T?�ӏ~�"�7j����$���)V�r��E��U�n�mA	2�����l��*�f����H�{zq�p�s���B+��co-윊��!���N���W�к=�H'R���ʨ`�;�ضU���F��u$ާ��[��c�y&C� �5��F}�BƸ�s��A�*�4#A�}4J��ϊ�= Y$�K}L� �WZ�����6%��x	�R���.K�i�Gp�
�s*estkN���pЛr�/$��,��8����c�yd���E�֓����.Q�7�	��yV���%�"'�ז4�Z)�E���b?�t!]�[�6� 	����\��۰� -����˷��U�@ƺ�����r�70s�r�3��dVRE~C
�٥yD�+
˃��%�$��0�İ�6��ۈ����:��|��h1�W�m[N��N�-y��� ��ا���uX��`�-�H�hW�c�:����I� �0X����}���{$�\R��/]�/Nܧ��Q�5*�c`�FYw��s��cN�u�� �q�ob�sa����A7�5����ч�ԝ��f~$7U@~R�S��h�I�ǯ|[њ���=Ő�.�	��o��%Ǿ��l� 
�`R�00�G��u�uG�;�`�?)fE�\_Y���5�,���q
Wj�&A�/����?��c�L3���h����W�J7EX�2�[�#�_-�]���%�86?�g��r����>e$�U��!������ύ1r�l��|'���br2͞׈\j[b6�w9b�t��ϡ=LLsm7կ��n2����E8Y-�) �������2���6P���C��\����$H��;�����!ly�5��P����сY��@ߍL�:��6��/�Lۨ�vl�p7lq�J��l��+��>���M� &������׉��*�gK��8�ŁX��d3�����
�Xbg�i%��% ��0�`�0���k|�4�No�ɏt��Vx� ǽ�����W�͎�h�>B�2�v����X;#WXmﲜ�tc� @]+����̮�獴i�~�dK�8��o��9"�k�m�ic���z��ZgO\�ʍP�v�����Qy�D�Δ=��b��U�q�c���m�����o�"�Z�ҩ)F׻?��j�3��B3SB@"��5m^,d������y^����>��9�����c�Q�|��X��R=7�ԑ�"t+w�9c�_��=�sԱ�<���XƘ�ͼrZ*�	��nh-�B^�ܤX<\�n�.�;Z()x���%~�x2��_�h���W�π�{=���6�l�X��Ͷ����Ȕ�=�'j5�6 ���/f���Ag���\#԰4��TM)����ǐ��Z�@���g�ki�d�ƺ�"������gԊ��6����?; �}����3��u晖[/
�4T�%�x7�5��/b%�R}"�j�8̔���`�j��J�����<�n�:��y��H(ڲ�:�x.��fL=�<����Pf�2�/_$�a�:���[ey���>�;X�Me�1��.�M�3��'�D������b�Hp.oG ��O�m4J���u5�b/]�.pg*	���Sp�0X��O�hָ��3~��i���*T��@|}�a�Y�q.�ӸĴ�.Ea%�<��	�B(xEr#� �G<��e=�߫� p�w��Op��e�T(����/0O��	�Tƃc��Z�u���p�)輷�.�G3��hࡎ(=�?�0OP�%���xuD��-A�FB���LL*�~d_�ԫ���l��(��6�E3�L)B)a-�,X�3��F�d�o��?~dYjQ)W<˧���fő������+�h�3&}��na8aר��lO�<�{��;"y�Q�j@�ݞ��{�g�puыCZA\rMϜ��ר���,�}n�S����JXP8o��H}��>�q���q89�k��o�2��=�^�\���w��#>hH��pVc4�rl�݀A}�Tɵ��@�oR4���&��+���.Lؐ��ͥ���Y�{4>����g�Ï�o�Ҝ�w�_2���@?� ���Cې|`|�����X�t���!9�5�6\j���I�i/�_7()*� 2����/O�ޝ6?u�!	LhGj�D�;�&�bʱ�����B����3���A�)i{-9p)g�!�?:����۞�DC!Y���]/4������P)\��?�5:�֞�,$S�no8�g�?:��P���X�8��!ia�>�����'�	��f��4|1m尝����ŎW�5o��O]"�����r*5�f
l�*M(�ARf~S�2��.yd�����28֏�_�n��>�*L��?R�����d��B/��1R�gb��lwu/��E�7�}6%|6k��M��a��}VYn��u@ql��P?���2:�!W����ð�4�@爙a}����^��G�}��l��2���)�&��3=�<�䗰i1����"H�k=c��wF8r�F-@����m<�������;�{,n2�9q�]���9
�=bD(�*��%�PԎ�n:B�nk�A�%�OU�g'>�g�[�g?$x�s�e)�]z�����%R��J�E�蔈�k��xB�?A��
�TCbnx�� ��ލ�H"^�<�(��z�;���$_4͈�xSӋϮ߮���`*������~e�EJ��p�����������	8�(Y7}���eM��J�s�O���k�#�"z�n.*��T���)UGz�`�m5�i��j�a����`����X�tI��h��Or_o�����`��"����ĩd���~��TOr\(�������KY���Z����+�P�k��o�a�Q'����;�Uw�_����-�#NJv.�Na���3��Asf0��0oȫ�Eq������Z�(�w�\>��냹6��4-a��C5�ñ��xUi��dhR��>�B��
$��$x�Z7��\��1A��Ȥ��N흿j� �D$z9�o�hwx�4��L<~�\&��� ���[T�g����锽�y�W�s.쿽,b��(��虥���zr�K����y�X��)_�|^�"1��5����c�4�<����~�����n����T�b=ųw��������7�;��4DV�'^5�{���
1*%���}��I�,����ҵ9�(U��D\��	�E�2�r'�	J(f�����kŢ�c��x�ۆ���0���-`0����v��kY6�/T�q�u�8;�NQ}�gcM%4}����?^���/�ݨ�I��a�鼍�ZY(�d���$�+~��ݙ|r��(.s0�W����+#0�cPz�b��\�Lw�]����{��2�����G��ny�C:�t&�+T\�ȡr�F���1<�ЭXjx2�����V��?M��%?k�� �Y{[C�d�+S�r��|����r� gO� $.���.
�������Qhr��Xq�|��pUS��:� _jD-��5硡�rٝM��j�Vf��/b�t�`�xr��S��ڜw�^W+M��pbkSA��E�6���\�.��EY_��R�˷���l������x�B�!�b�sSW��9ʬ�i��b>�Z�i8���V�y���0+[������óI]X'*$ZS{�{T3q��ALbG�nAC�)�W�M���s��)�x���8Hoiҽ8���2]��׃�z<zP�?>\S�Q�ʅ�qדl��r@�(J�"���2$�]��w�� �3�7,E��[PԄ^��'� f��I�b�J�<lU"��.�Y��q.��T|Y�?�%27'T��Z��n���?c3�ĬX�o~��H�����݂�x��s�\���l���z�K���a����~�$�i���7?ߓ;\�F��3��-�'�4�^�C��\����Nс�_����hU���"�?�0���g/hf�'�K$�X.dp�-��@_}�]c<��z�L}8��l�(~J^�
���cE+��1;e�����7�z��`^4a�1���OP(0:�	%�:;�q�W8�κ?Ul#\�xKb�R<��n��^r��fl2���db��*Lf����
�1h@�i
�S������"w���pZ=,�GG$�ŻFh�ۋZr�� ���`: ��K��/��h����U&^�Z�b�����h�����d�������4���}gn��@�����.���q$g�9�1�������;��(ia����`�U�b�W�^a��['ݓ�&���wQ7�q���?.;�Nc+b}�h�T�0^�o�<�a ��CX�r��Z�� ��6��Ĕ"֯E<�w퐪 �"�F��^�s�M��^ҞErk�N.��C��|f�&�d�8M{�:!�<-t�4j��ܤ�\}{0��j��m��u�ЅZDI���\��U���\(�1Y��Y�f���;g&���U.jH]�����哙O�b?���+/���[�8�,�f�X��D
_�*g}��!�2S[�S��S]�G����lo�(���0�����k�f�j<lV�э94p��$[�w)&D�
,"��9�@7��<j��?�2��Ƚ���6S�sG$��a�B��(�|���� \y^\�����%�:�nY�U��Zʇ$�kg�3�!��-� eU }�9���fo�I/,3�h&�YFd8��R��
���a��dي�����S���\�����3������߼�Ic��z� �8_\Rڷ�@�l>����ҷVw���H�, �>!N��I,/1������9.��-���U�!�-�d�Q`�6_�}��!b���! {�/�P�Z�2M����o��@e>8f�aQڙ��O0�W �D����7Ȫ��D�$RU����AD�0��H{��2�+�Q��"P��=̀����t�����b��Zh݊��~�%�j�������F�%t֑���]/�����{��:�"�a���@��1�X���N�f䎜T+���+
��+�Q��������:��2��;�����'�<	�}
�7��q�����k�*&�Q��h�t���
}��c'/��O��#G���p�`2,�\���V�]�]^��� ��ȆwΧ�J!W�$j�k�����[�3U�v�f�����Ȋf�a<�R^�I�-��At�Y�P,>ȌLw��$��.�Jz��X�E��Z� dD���#�o[k��3�p�B)!Y�KAʣ�W�&���0�q1�r�.���ׄ��S�@s��M�c ��� <�S݂ל��~���+}�Ns�Ĉ��1>$���q���g�sM���3�D�!��`��m��O+�)�Eď@�f�����Tb:�a�5��=���I#.Cʕ��چ���=�~Ӊ�z.����ao��,&�ÑV}�p<@\v�<��ƀ���ѧ�k ,�N"DnSs[������H�=�A:t?^�i�v`���7?zPP��IrCI��RG�ϸ���f���q�����+�3%f��㯮���"�p��[�X�2�WfcK1�C�e��Og�5��՗I�P���h��R8�?c�����9&5U�m8�,ԩ��j��>�<�|51jx5�T�F�?����2�"�� %]3W�N%��,[Lp>�Y��=	8���PG>4�g��҇L*]G�;��fP�F��9�b�B�"6>#Pmmxѕ�U��FA1��MȂ���hC���9�ZQ��q^+y~�<�ue]P�����-b@�|��vu��T�b֬^Md����ӹ���gW�̻�t�=R��o2��eSo��u�A�:��L�DaGn�K	@��:)��crJ->V�	�F4��5䷟h�o��V�^���	�!���e��NwZ�H]6���QW&XV4�evf����
�&k7'x��2Q%�d�ːEm O_�=�؞�g���OBT���/aXs4�h�m�o������]F3�
7d�}��p����^y�I�ۨ�#�vUZuj�d�ИFO�q������%"O�jHO����=�v{<m�7BM����U�e�;�5�W�V$��������
tde��H�1�Sqxᥪ	������)U�c�Z���U*8��J�)$̈j4׃K����a�>�)&��=��_�vF<C�joC]ͷ�l����� ~-��`MhP7�6
3�\Ϣ�dg7����b�j(�g[_B'��#���r��;����\�D��ʾY�g�9-M���7)�8�ݬm���;��U�(���a��iu����g�եKO��xV'� ��vbn]+�ħ�����髭����R����H�un��Y�.�NlY�,lI]�θ�+ru=��۟y9M�	���"rˎZ�f�S�J3k�'�'�k|���DJߑ�J�y�>�~�ǋ ⟵�g�R��-vW�н��,�p��jAĴ>덙v���5+��R��Rc����x�da*�8ۗ8�;�9��a�-��@��Y��k�Մ�Vwƛ�)-F�ȑ���?�vp���6&�:�'h^��v�D}0���B��ћ��8FQՉ����js�c�=������?/�O�����l�Se�!��'�H��[�(��@XD�-/�_I˃Z��<�/�z[n��yCD�@i��D�5Z�s���r} ��#�?������nnנ�NL2�lɼ��9���5xO��� oL�A�jt8�_0V3t52����eG:7zF4T�m�O�+ǚ��,�5w�}�wX�9�`ݟ4N�*w2/�Bǉ}mp�Z����	Ax˅k��]�e�V�w�Q���h�&�b"�&�3���;U�IA���)��%-�F{ɛTK�%��܈8�;Cn9�4�rw*�����ː�09�D�������^rp�.\�"�{,�ϓ|Hu_#�x����ښ_��l1c+?�R)YYaD�?1Ej�w܃�i�=;Ve�Ue��H�jgn�.��
|��dX��h�	L��p1r�n�l�De��}	�bJyxw�j ĺ4�9(�U)��,u���k�ܚk�L�����d�p��aA|໌��}<V��/�c��VW��{�^C{��[we��=d��V))+F ���I *�1�W�4
~<~�4ت�xl�KP�W#+1|�W���J��o(����_`V��y.��A�,*t����p��A&#a�1y��;�g!TQ���/X��+D`x\|�c�#f+ۈ�b�f�F�)�f��:qt�+�{�5eq�о��{l���]���x��a{��ѳ;����`���;�ց�?���#AU)(���*�$�W�v����t�,s��%	�y��޵�*�Q��DR�-���6=&�Fb(��@�<�����MC�x�zO֍��Q�W��_�N�a#A�e|S��C�m�~B"�8�55���	|'��`�	����)ݘ9�Ŗ9��J˚�/�����}IjʥL�Y�~p�(R��,�*�ͬ�O��9�R�\,��- �5;����*k�e�{�ߎ�9K��{��<%���R�¢<S)dW|�t��w��Xt!�����4E��.�c��Ӆd�y�B���Z�0�Ǟ^X��A���H_8t^�$8 څx���f���?�#���Fh��^e}B���M:e3.4���pP! S'�=�/��X���F��2��u��;睉
���8x�鿃��;�u*�T��g�{Ȯ�	,���3 oVͶlv Ũ~�#y�ֿH��｡%~z�x�#`n5'����ƛYO|,ӽUZ���BpJ+��fF'��Ά]�z/�d�n`�,T.ˮ'��E�>C�bn'��TPv<R��5��o��qj�DnG���pVO�'�ͬ���f�����&	 e@��U�O���OCU|����%�Đ�Q_(@�.^��ہ �ܚ��R�:(S<��F��;���a �KD�z9,��2�h���s���s�Y6
�㐌j���"����_�[G։|c��1D�
�����+���֐�Y\��'���3�
X�� P��줣R~�~dW���n���	����J��P��u<�)��
*�zr8����ᓛR�Y��O[b���"�먎|JnD��)De��zM\*��6 Ok�Q�'�h�sm�v�}d2��D�qFx���#T�!�:���������,�=���H���S�X�E̓؄i����f����=�ŗ��՝������W#Q�BFۈ���ŉ�7ʧU�'�c9N���+7�G�s16t`WeqNܑ�����ti��p���a%x��B�d/�xʤ��
�P6˭x�I��@	�c��.�}Awo��(,�+۱6*f�F;W�΀+�H�>^�m�S�]Ň56MLE��2���_g���ʁ��V�.��V��F!�o5L����O��A��"ֆ;�_
@���dm� %��)��Lge����#��s�/�teNCT���:,�BmN�~��8�A��d�g�`.
��.�@v57����"��|G|���C	
��rn@���j�C��An�5(�k�	��9���n��b�,z���x"��Ul�Ox��<|�7��^��倍C��-btm��$��0IE>_}�F�w�e����q?�$V�<v��N��w��:�������k'}=��{��hc���x[ �&Oi��Ɔ�j���^`�hҡM�k���G2և�L��Az���/���Hur6=6�vf����Cv"��:��u�f���`�|0G�4�?��K75�"����H�65��Z��x���f�	��Ǭ�x�CJ\�Ƚ��
�o��(���"�݋��޾���@���?�3+�/�+� m���&1����4H��j���|�͙���l�֊����S�����ᦲ����D������[�%՘|�U^�0���D�'ˠ����UN6�N����t��@���Db���:���@>�j�njp�d��Z�(�R���%֒Y�w���*z��-F�1P��an/a�6�p��1� �_�y��%��'s�%�]8v��D�ž��*�d�5�nL>��F$$cb�( F����$��L���R�R]�.]I,Ԙ ��ϫ�a`���K*�J:#n����N����Z2����:8�������/��A0e��qE��C�.�=�Nc�)�{,ܪa{y=L����N�Gw	'o�ܘ���a$��0zit������c� �&��F������O��WBH�}��V�s=���g�2CQ-�E�Ԯ�ح@���6�:b^v���ZK'�l��<��%��`�D>�~��v��C4&IY��*�b*r� �&.���*iO�k_���^�y,�~>d�P/��vL��tX�n����]5�8��>=i%�d��NBr� �~>����w����T���@�~p_yuw�y�gi�x�և��R
���k��滲Y���fFteP�[s��0�/����AWtM���V�)�M����&0�L�:��$���ѕ4�W"��Iw0) B�'�սd���� ����L���4�ּ�T���ο��IN�;!>%T�ER�J:-���cV+�j��i.�f�C��W5�2=�ʰ�P�>گY����o��=y�5묲�b��ҽ�'�w5zF�-{(��Gy����_9�~ڲ��Ȩ�j�O�qW�a��}¾I����r��`�7c�>��%��a]*Z�[S�� o���և���ͪ��9�P1R^��}��!�~��������g�=a ʦ�(�EMe������p�C�~��^����T;v���!�p��ǀ��+�a�O�P��̫�{���-hS����$��dһ��ǎ=S��h�Д|;Ig�������ln:�*���v�rc4����&Bz���c�������3fj�{�n�?.�sD˰<o^I>3-�h+�C4ȣ���ce)�A@2a��!�W\Ͱ���/4�w��>�:ꆫ���[֊5�	�����n�z�ã���}LW�]5�|�R!���l'�x>���N��4":q�6�Z&��a��*9;�O%�v�3c��t�+&Y���$g)n�������f�*$�;]t�Z���d��/�	G�Y�ݍB��Hn�4ZTC�ӏtRIF�o�g�e�R�_z��3ѸK�P�nW�/��-#�Ɏ� @F���"���b�Mv�����:M��&������-	GO�>�e#v�>r\������lNK�a��?����O�*P�S�^�7�OT�r2w���J���ɯm����O�H��{�.�d����%�4<��psJ����
�\�h�b�����leB�Vx�d�J������0�jF������tfޚ"[���a���F2f����M��[L��;��R
3JRj�9�a�?�7��p�n�A�V�H��$=��@I�|�b;�V3���`�(��\;�F�աw*��[�lA�w�n��rg��|8K���(�-��}�7��vQ�3G4�_QztD�rO�BwvI�k�R�'����W04B���3��� ɸ$��?O �H�%��=x������oD�[���3�|[�0�v}�riI��v�����e�R�\aw�\�N�~��a$��q�hi��0�N�)��7 $I2�K��ͩڨ�(s���t	�7�)�<"�n��N�z������M��<�v��W"'&�5&� g�� @���|���n�;^��*;��E��8��h�P0�Œ�tob��/t�y���K�x�2-v��
�!���eG�:�;��̽W>�1k^_dO�ؙ��LFi��x�"!�����ԝ�v���M>�V�-��U�G��ʑ�'����>���,;�q;��<ċ�R�~d"���'^9d:]�����Й�r�.�z��y?[�~��h�5!U���o�&1���m�`��nG�{�~�{����#N��g�Ge'I�fѨ��� IY��b8��\��t�ne��&Dĉ�6=�%ɏ���~о�ze�Co-�_�T\Q*��
	�a�.�B�������}@{��e'�<~c��R�~�S)��_��>u~��o#O����k��y70�Ǿ�0����>ۨ'(iLV9�H����_�:'����#Lmi���/�L�2ir�o�_���K���ǖ@#�YN�L��ES���
I'F�uE\c�y $<������i��s���AD�Nn�D,vԌ|���� ��8���y�ԡ��c̍���������n�z7�M/��0���AJ�7���?�}��Ɨ�8GZ�ux��Xi�+/X��g�w>����Dx>����A�L�[i���<���V߰o���gK|���,Ol$:'�&�����"��v�,�I62�Ǩ4���2����ǥ���!�ta&��g�N\0p>N&c����&�1$n �V&'ùam按A��e�J+�e���&Ag#�%�6o���m�PA�;R�3߶�!���ޟUo���T%U��1����FzĆ��kE-�w+h�G �O�wXI�y�d����N"�o�f���_z#ܒ�^��Ր:٩P���eQ�2���a�$�N����^��^�P��!p���k�Y*#�8��Ύ�`�ǻV����F���Mg��B����_�k�ڈ�-�&�iAr�ⲹ��I�ĉ*6������GS��Q
NŊ�����H��p�F(cg�2�8͌-�n7s;�:8O�bc�S��VC�mj��5�O1���2��mq�1av�>����Lm,(9E�I�Q��G�9�PW����&�H�4�B�W�.����
�f7&��!�\vnr����#Y����:H���@�;�A.�`l��~h~�|��'F ��
���g:�H��Q�<�O9s�'�}�4�pU'��e7[�)�z8���)&]sE�z<��C���WVy�.��:UN�k�Ȼsҍ��M�����)&�]_���������Ͼ[��nU��*w9��qU��
�J�5~�Ⲟ��y$�]��s(��!l�[����q�c��̭*RU��p�I���mN�{�"f�?�b�r��25	{��s����nN��y �
����]��'@R��ߠY��{g5�w� �1���f.wV�����[�BOr��������s���H!觩A����\R�k�P�@��~�]�g���A���Lz�?_�|j���#�Osjh��^*w�d�ÖcA�E�FM@�����7�g�ut�n0��
����b����j����-E� �ѓA��zG£a�-!���v��V��u��@.��ԛ���`����]�R�
+�2T3�B�,2�0	����������bs[CX�VoeFp5�\�X�h3����l%�aΖ��ǰY��5y)�k,k-�G���|3�=ﰻ0rj����pk�bpn�)�pE�K{z%���(�����7�mx~���i��@/��g'�Z�a��®��J��8�ٟz>[���E�,ȟ��=5z
v��kRA����M� p!JW��8�8��D�lH�kP��_+����~��֩9�3(��Jv�<s����e�%��ݐF�bE�����l����'�@�7�:�L{<�b6Q��!�F�9��a�)�jߣB�l(���ǎ��>��)���/5���H{m�����w�	p�����}�
��K\@���<H��<��9.��A��G\t�;S����w��r={Hr}jB d*9�`��iIO徨��pR9i:3	0v�{@�\7x��U;�P�B~���F�����WVXw ���s_��CE�ډ�_3���J{��D��de'�v�ɖeန ������0"�oʚe��	ۨ�����')}Zs���5�v�ܷ�s��}}��J��6���ر=�{�._|��z�k��Q=�櫂|A�*zB�������_�9�O&���� �2
������%�S,�mA�X��QC"	 X�?�����\����Z�-��ֲ9�S�:�N��(�1ѻc��Y�p����"Htyo:�� ��dsC��90��X/o0Z�h��RT���l# �sc�a��1����EX�1�p_Qi���~�X��g�0!���L���W��lw��|t�����Po���L�-���h����&��Cg
�"u�eY���v�82}Z��i�5�P-�ꤱ.9�05F&��@�EPC��n�vF<�̆��ա"L�˕Ʀ�i�a�~�?�e𩊾I8���	[$[�n���Q�d�1��k�n�n�4��ù���-��O��^&{��wu�l0��Y�4����G���R�SSӟ)A�瀝ꡄ����䘙�����}�
)�7-�"�	�@�	/ggv�@�Ag
��zg͂�0W.�����q�8ԗ���ҎbTm�;u	ˌ����骐�Qѐ��ZCo6��)��s�pw7����Q��6g�%jp&�q��_�EEg������G+2�BR�H�7��,�����G�0J�x��ʑ��	�ւ��{:wm짋��H���G��9p�\�vco���X�.0���%ޑR5)P���-�K`���q,SſEO���5.�'�Y�y���Iх��O����B���O�$[��6��8�6䥸�ERvi0�p'�[G*��2P s�=��V��LH2(IҰYD3?��Qo�~�"(� ���zM�^f�e�_�%{':xY���P���,�U;ΉNsf���Vٟ���@�΄��;�Y�\a&�!Lwb�ur	��r����jw�z�K��軁ѫ�3��ȱ��i|�5?��4�^���/L�M���eV��1D�O~ ������<�`��n/�A�% ��څ��tp��i&3�{� � �S���_�\O�;.s�S��;.�oJ�HӮ<�ô⦳pe�'hA-�yY7�͞�#$��q[���'�Ψ�@�y
�0���Ef1WֺCu�qu�*��1�.rې��<�p�����j:��A�:���lܯ��|�M�p�D�Fh'��&�ԃ7�;a-a�(8�DD�R�.�,x�����Duy��q���K�_��	���#�*���j���5\5��<�c��+f���չ�����?����7R=
���3X�<����Qz��o���샂��J �''݈il�	��<�q��W��A�I��m�~r��'_��I�S�\�L�q\��A76h5U��x��Ɇ��u�E�c���߃d[��'�+'@�n�F�ۯ�ga��ɚ!�uЉ�;��P��
%Ò��65>���k{u�ŵ񙞧��aְ�"̭����%G.Ҫ2���R�v3_���Z����1������G�åln�� �j�r�8
2�O��FC���,�7f��n�VB���"/Maˣ�O�se�B�Șc�돩���͕G�m��ֲ�5�e�y���=����u��2�r"��_0Z���}8-�
ղ��<2����LȠ�=W9[Cj}'�m�k���LIlHa�ӌ����*�0H�k����zL��K$�H�U��Z��k�=+\B�{p��9���U�'#8N���1jC��F���Ec�M��F�x�j��l��fI�5��h_aJ�&�.Gq�id��uð���s'-w�w�=�T0�N��e+�C�焓L�~����k m�;�ő�ꩢ)�'rW�;go.w���R�m����'�a\�(���C��>8�;C<��t6a,
w%�rzL����b7�u&����f�_�����Ig :Ψ)��33Qm�K-����B���#{'6�vB��R�0���лg�W��D�d������`�nm�-��	MV)Ut<$N���G)�3o.�����"��!~DP#"���=@�|�mV�6���߃D׭��2eD�)v��lO��6S���j:p�P���{��������� +?Ԣ�M�,��(VFׯǹp�?��L�0��#�.�p�	��p^��T����8���i�?�Ċ9%
cA�T��`�Wc�ԓ������[��3��^�-��7V��%g���p G��@�O�j�*�Aq�Z��ve:b�2G���d�9�2��=7N������/k ��b��-8	_|h�����Z��ªR��4]��#QU�2�ax�=�$.',���F�`Nv5�v0Ic���.��t���!9�7)�zFA�������gI�,�H?͹@N��>���юU���8 #<{0�A�P9�s��=S��?Lw!�n�Jp�z��E�5B��}�3�w͙��6��7��r堉�����[PJ��yk+�D3�-`�+�g,N�	jEb�k�c�q?�5���+���i6�F����Ë�B�e�a������J��s���t�3��
ᑱ���4���BR'r���j��)S�M���ℜ��X��;Ұ}ʓ�f��^K8:L��S;��l��;���B�䊠��l��Ϟ�]B{������T5�Bt�g�X/u%��&R�\b�*��+Uj���$BE���4N��.��r6F��M��;)w�������ye��I'����l�I���d�"���w?��y�:8���&yE+̘f���\��>2U9�t�`��F�}�k�	z�k3fkbK݁i4�8k�I�Y����@X5K�.����m�_#g�U�o�ySˮݳ�-�(�Akđcԃ%��i�����.,?H��=�����]_�J1B��&�R>�_�d�Z�3��R�!Ǔ �C����R�q�����k�������9p��w��%�DBcv��$���f�/ӼHs�b��#�M��L�D�^bG��Co?>�ճ�1P�����p}X�=ɍf�<� >���a����s0�E���kNotqGᯋɏ.'x9��ۊa����+@O�{n#pu�7J�Z]
��4?D��O!x�}o[�vQ��FrzOU�o}�Y�b���i�%�%�yl�b��̿�H
�y�=3^E)�*P��/P�ys!u�v�;�}D �C�w�qbt���^�i���^ǎ�G��|�#��Io�Щ*���Ǧ��ވ[��j��Z!�
�W T�a����6�+zJ�<%�r��=�ѵhko�|Y���k�K�_���@:�1^T��c�-�26���{܏ [e�q��C�Ni�9��|^!�6�����9��)���F�ws��nXg$v��T�����<�Sh���DMg�6AP	�w��C���Ij�{����j�[��_�`��@��¡UHܫ-��G������aLXaEU�:]P���N���O���e�%C]�V{��-1��q9�<X2K���[�t�t�)Bϝ�_v�v�٬��=�%}X�pœ���r5J�7�j���7��B������9�.r�m���V>��`���X�4�u��v�Y��)tY�u�E����	ɩ�,̙>�3��wyh��}G��X��~A�;��_�n@<�B����;W:��v�!V��`�kU����+�yI��ha� ��AE��s;�ٞyJ�QM��{�4�fq�>�C�t	�0�!�"�;A���@GT����'$X
V!m�O	L<1��.<����67+M�q�����
w?_��16��y�8	!l6�X���PH� �'�L37g��!Y�1S���=jCP��(,����͜Nh��*B6���hs�y⊌��9�E��)MX�7F�j �.͵���! �mh�񣜴ߚ�UyI4�U��J���f��a��K�w>����������}LݺJka��`^�_�q7�(b��1��5�������nZ�9,�ڪ��M�0��J�aOsp�._@��+B|D�����S���'���Ms��'�����i͂�nG��S��Ԏɭ7mNB��sݺ��ܾ�%9k�� t��:��vy��m��vJp��~XfぷJ��4�cDMT�S�KcWqd��)�q�+�Mg�<z�������i�7�Pӥ8��rzD�{�qvh$ťw�L$"�ӭ�W������e�f�ʋ����n��+�%m�0R{���;��S�͝����^��؊ h%�C�i��Q�1���l�;5���eb�A���U�8����D)E�OxGln�ڤ���E��GZpz�AN�瘯㥼��F
!��6�{̩��M�5��\"�J��wo	D��E�+���q�iN�O�绡������72@/�w���u�`w5%'���MU2�'I9�'�}����>i�W��b����CS�G ̵�\��ƾ�m?n�7~u���%]��,)�_g��_}l·���+��e���I�K�H)����ZLu��Gg6�#�l�2+g&�cdY0�X��I�$a�ZYU��T� ����~0aA���`-if�Bg��7Ii��<[���/Xވ#lB��*l���6ۯ�bl ��ծ���"[n�+��(�\��tY?�BJȰC�Pqu�a�PT�p>R�
��7�+�۞�T0��>�C����+T�$�Մ�HPy'�0�)�
-�a��`��=׿�y�#H�Fw��9��]�����[%�-U#z�1��<�H��s�G�_�e6h��q�)�c����$S����9!Z�~ H�sI�!���uy������e ��V@�W�zg���Bv��D�=��Ir�<I����6��`D�p�Ǹ\d�������n�6��w�c�3^L?�
o�;�e:ִD��=32��s�An�r�f:n����I���xb��cZwy3��H�u��h1��9y4[��I礢[D��'���yEL43�F�����#�����l���ʐ�h��.}�L��[z��ǯc�u�S5��{�u�@��Yi�~H���4VF+�����sp�^��>���ۼ������,aog� �7�T  #?�䯦������BC'��G~"�q�[��p�lF�8>(�����q� pVБn��MC.s��6<��.�a����>f<�]���
�\=$^Ffސ�0�E�!]`�o��ϙ��pc�]QuЦ,�D'��ro�jh��#\�xu#���(��*�
	��Ž*�kv;��ܳ_�|W���s����S�>����J�!����>�i��?�*#��p�~��6ɍ��yk��b�ޅ�4Ӑ!7�N��g��X��E���~��Ө2�;�k	B�*c?��}�� ר���4��F	����7���\
+n��r�?�2��~�J���z��B��AohXB��˭
e(� _҅Sꦞe�z�!�&�8=FjVO�;绒P��|���{Hױ��3��l!�$"�<o3� �ck���REΗ�1�b� '#Q%���<ms�yՐ��Y�|E��5 �v�n�
�Cx�����+&�zf�Ea7k�'�~���cJ��m�1�<_�ȇ,՚��t��=��
��㉩e?��=Rg�-��R�'e��{8m��WC�=<�m�rT�P�WH��y�Q�2�]��y"���w;t�Q�q��܂_�Gi8C��n�~�#�s��}&ð���ºe;���>�F2��~|�q�@�5U���v_��Z@$m2�H/�l��iGF�Y����ēK�����ys�
0��Y�	$d��[�K,\s�E@���L=�/�ڍ"�@!���0���>HZ@�^�!L��J��j�L�{�睃ŜMGL�F�唐��y%�:���S����W7q�C����Ψ�ы:��̜�3�K��U�-[�^��Ll�;���2�9%rϳ�S���<���s}
&{}V�y~���*��c�
���*�u��ա��N'zJ�Ѝ��=��V�J�R�,��%��0 ����	��u�b�2�o\��[�%o�us<��=�����d{v �d+�+#����2;*f��<p*ROJ�#W�A�/w_ѱ���@Y>q�;P[^�D7�; añXB�G�o��Ԏ.�D�҂�9q�J2;�2VjV*g���3��/���*_��G�M��p��6��C@�l�u��]���O���B��n�zl�S�l͆8�t�ۺL#�}ńZ��oE0��x���j!"�_�P�
�;u �C�_o4: ��24)�`c� �QI����8�@��[#}�d��L!!V�>Ȋ�p[��i�la�/k
�T���b���1O��4%��N�=�_3�����B�f�ѝx�28���а�=˰F��IڧͥB�k.����S�ފ"p����C%W�&�Ϧ򁃔SF�<tN^�����ϩt�����M�!��������]D�Gq�$���v�P�څ��p���B���	%���'@�5f������ X���w�u�{>���S37�����q��[v}�����j*w��5�5�a���<�8�ϩ�:�RF����b��ö	L.>��P���Z-���:&�E-Ϥ�k\Ch�4���s�<��\gA��k�n�Z��v~��΃C~ׇ/����kzE�
��^�3���9e14����̺�a'��mK$��b��Sh[2���(-Y�׾>�1���t��Rk�����q�+}LDj#�i*JN���u���T��g���6B���B��J�7�=����s�g�[��{�h��H��-d�p)@�I�B��,D��sͿ.�qyn�c��\���iߊ��z�O��݅�E:
���Q`���Z�y3�1/|#@uZk+P@��P"2:�]��m�l�����)�Ac�q�3�P�pp���D�o]]���J�?ض��E��D����r?=�T�j����Y��y�z���H�;�2��`��KA��x�ߍO�ER A{7M���~m
r�(&c�t�;�(7�o%l�wR1�wֽ�}7	#��n���;�N�\V�,ד�wv1�����ju�j���!0CN��VEq�9Q̪8�[����
G���[\���d*��y��(lS1[аd*�s?ܛb�G!��o�v�f������~!���RY(4�;i䓐:0�@m�E0<p�~��\���*�������h�3�P]�b���KuЀ�t���~R�D�-�;��7(����V�n,Ӧ�6ĥ����x�R�{Fѽ�6�XA���e_�<p� a�����+��h��>�9�on����=��A:KE�SO`����ӎ�)��k���W��m��ztVHM#�-���5$	v$����X���q<��-|����CC���b�\�Z����qw+��9NX��"�s��gO ;�Q'ڪ_?�즴���0Lp&e0៙)�sA=)	 �l��	��z�O�=`Q�v-7��%VFxO��Kv�����Iɬ�%?�Z�r��|��Я���N�>4���?m�EJ�S蠛��Lse(fEL�w��vfr�<|�,HjS9ӄ�+����_�S��K� ��"�ӯ%�0�y�ɺ��Q�(��;)$��^���&�]�����-5����n��8�YY`*���F�G.���+����ٓ*)����z��Tw���� "�H�s+ScD��'�h��;�gtX���"v*C�����)E��Nn�K<��S!�{P:p"�)�lW�N=$-�y>a�g�4]�F�M������4����.��\�;Ub=�}�q����Fw0����l�mu���>����傝���!v�ʀ�w��0z%��K�q{E���}�A�J�M����rL�a�*�jB�=W�r)��������z2O�)�'�W	��A���%ym2�C�s:es�4�QW��k'��܋ Y��e�O}��Y����ze�C�%���/j�e ��B��L�<.s^'/�	K��a�/y�%
�Mj�R��[�Q$$�-��gf^�DXa~��a5�R�&�=�����������Q�Q89��b1>G�'�>0�ת�wn\S�D�[iss���4\`�(��fO������<�G'���!��9�8 X����?�u�>��h�w;e
�{�T-]�Rj�1GvS�=��.(Hi}���s|���|��7`D�����1���cz"�G�����H�NՔ���P�ĳUW9���� �R�Ὡ��B�d7T�#��휨�UO�#L��C�;h^�9O�{1y��\,�&>�	mms�o�h:����砠{�)��;Ys�@�Ś	��x��t��qA{��*j7�5��DS�����;:>$�"$W+���&f23����Z�~�N�ȦUܩe��c��(�&yaL8=��9�)=&`L�� �e�T!?Q��.ė{��.��D,
��$t6N��A$�y�����;���v�j�D0���`������;����KC��Ju�0ܑ�qV5ڸ%/"i��.l�d ��-�ɌU��l���@a7t�U���Տ7{ ��4����Y�` []�su%I���If�з��J�����V
_��wI~�j��;�h[\T�؇�L�G�=��0O耵4�������i[�j���z���s�S���#\V�H���t	�j)��R25��r�}q�
�iA�������$��hT2[��iN��p�ͱ�	�f&�Ǜ˲%1}`Ue�^�4Б��q4\Iq0��崅�#h��W*�.�����0��K-����>{(p^��p,c̢�Y�,�e��D:�^����?Ň1�T������4��Z���vD�7��c��aX��N�N33��K�2#��]J�� Ie�kYFZZT��++X���T�t<��G!YL�Ș�߶VȐN��*:Q,fwf�Z��0x�D��[:�s-(�!pX�w��j�?��v�7�!�,�;��Y�3����?k+���v�}�;��Q�G��u<W����C��+���2�5�ӄ(f�W������	�\��!�)��7�YB����y�n�@�k1*��%�@�V�Uס�D�<9�ӗ�26��[�vJݵ~��=�F~	t&����c�T/!����� @������#�B�u��e�b==�����kT8YۿGU�m���jPq��>O��Y;�(�~/��G�{��@�����$r�.:����W��BN���fA�_��gR� `���|���g�qnB���1�\���!{4����<KP�>p�(�1>�Ԫ+3��H;K�7�}�Jz�ڨ;�~6�cڧe}�E�x�{|���BpT��4x��҅/���+��b�bJt������p���~>�Y�Z9�'��.�E�3����l��y�~A�����É^�Ν���3�	���8�z���M��a�,�ǵ�7�e��%�"�Ō��p,"m(#j�{<�h]�Ŗ	Zox�8�4R\�D��f�+�'u������Qc͘�I=��/r�u������UC�k�D����Z�_r�Bʖ]�d�Þ�=^��*z���j�k�VP��<D=� ��os�i�N�RlMA nG�[����<��t�����B�4i�Z)=ҜdZ"��ɼ�O�a��;�>��3�W:�8M�e&������RX"�(��LQ�;�� ��>�șp�ϟ��4���&�{X�:�4���n+�k��"��N�k"�i�$;�Wo�Ft/�Џ��ɉ<GA��b�1h-���ܬ�$�Q��2��ZM�ӭJr�ɀ�8���|A˟eu)�.���D���l�P����;��9뻜w��Q ����h1�n���l�:��pK�d�1t�T�����J#���b�����$� >{%$����F����&��mH�����,E�ǆ"7^������_D����9�A%}.Y���>̳c>�WP�"ᯞ���UL�����>�'��_�a)�A�����{�:­��m\j�ᷥ������5���;�ɚ�*�A��?|&4˧ԻN7���l��.Pߚ7+o��]�f�����P�p[�s<���T �N��%�bY>�4�U�-<i�H��gG��4<��t*�V�:	q���:xH�[���	N�>�۪�19B�u<>�E>��>��Bo`��4������1��iZё&���ͅ��%Te%��``�ϜE���L���|�D�\	�C�i��#����N�sRA���p.�/{h����"��KQ{�n�GGi�E`��TϚ�h�!S!�DHsA�z���b�c�9 \��H\��l@���U�]�Ee0�:7M�5C�{pZ@y,�5�1B�9��!R,���9�69*X�UC�ڞ\��n��3�ٷ�6���/3���H�ktf��"�h?Q���B��M]���.	$*K�͸	EסNY=�%���ߨv�"n��]n�L��JY�X;�9��؛���i/6�@}��Qdg�S]����>�Y�HݱeJ}��.q0�~��f~n$^4n��a��&��kg��N����SuL�i��z9�O�K���~U��f��Mz��8�
�y��҇�D�y�����6ػ�T�x	X����O�b������OA�<�罞9pZNJ����p�x����3"�Et�|)����6]�K�3<.z�J�?�{�e�,�kG�k��� ր�F%�J�Xo0�ᦸ#��}��t`����1���w��l�jd�n����E��v�w� og�@�$(�t�����Uc�P��^���oĥ@��/� yȊ���X����R,f�GQf�Ԣ��|l8�{��^11l��A�X}+|�K��0�P�:��I��>b,�o�~�e��3ڛ֢��u��Y�YX�>@m}zaT���a\}V�?S eD��~K�t_e&8z��c�~3e�p���d8#����a������K�Y�4O�'#���V�rɐT���sU��H�8�=�_�e��8˗>3V�0�A�!K@��"a��Q��6;i�4l�� :=�|勩ȴO)��d<JO����N�`�0(Z� ���q-��Ör0�)��&P�A��@+
P��f��޻*\�$�t�H��A�!�%j'�d
a�[�K�6b2EV~2V��)1�����l:,�_�NMcY8B\�G',_\̉���m��n8Y������C�q�7P#[3D���}�'p� �Tu��?���%G�S3U?$���-�#������u��nr&PsS��B��w6�"��]�A�R�!��Y��l2u�7�DH9�|��󳏵����K��7� \���
'��j���#��s>٩��W=�R��-���:Ħ�;ʳ;�\W�*�]�d�Q�l[�73����9�y�����1͓m����H����1K�r��K 6-zN� 	����;���(b�њ���Vu�I�Yy�ɠj_�W��6���_��;׆��ཹv2�n�
Uqݏ��󈬫qj=�V:#Xa�qZp|���5
�Zý�N8;
%9Ҷ6�$���f�Iw�<�����_,���9��N�����̦M�ߓ]��/39*����Kl���*�DsߓI%��p"K��޹=�#�B�H>���I2��)�Y�8�8��Bg�+�}@�&�p�.R�}�a�Bfg�Py3�(�{U��a݅U̿<B��e�L�o�P7�ɢS��Xxb���@"�T�f���
&�"s�r��N���4��<�*�3�� �sė�5��?\<}w��꺲y��Hy�ޝ�v��� Ҽ�q��R�/�c��3r�2҈"4��-?L��
F �� ʤVcā�[�e'��7�G��L^������ڈr��<[��?���:o����WϷ��3�ǅ��z:F* >�!��q����$�P�V(��F�4�Z�qje��B��2����a�
lb"��l��Y�å�(�`���P~��o�i�LD�XV�ΐuA�"�jϮ�ڄ"��{Ӄ�ۙ����#բZߺ��c���O1ˇ��9���8��V��M��(&3B4�ʘ..�� �懵�H��Q�����%S�k�z�U� �-ue��Aw<��(uJ3Z �YuN�=�?B���� ≋hM��k;��`e�'���w"O���F��C�Pv�ǽ[z�5���_�G���'�>r�"D��z|�T�z'v{��W���Z5?�q�Һ3=� wQK��z2�8�Ä��r6�����;gd�"z��NN'�2c�4����WJ>���҉����ܢτi�`��C��-	,�y&���-�9J٢���y;|2�|����=�+�(N� Ǭ�q,�����+��>n,DQ�#J؛�=��Tkbu��c����g�������K���x�F�`N�9��wD%\[�%i�lj�_�r7�?�]+��rC`#M��p@�(z�y)�˱�M*�:��s�ՙ�f+:�} ����4X�MCPV_os`�������tn��A�/$�־kq�sWΈ�&����?B^I/iN(���b��H�J.7ܜ/�>Τ;mH�~���>0'9jg�r�6:�P^�"tL'�C�&k�LU�b���:�QH��RwI/tU������>V$v�	���:�ͽdNA:H�n]�d�~�S�t{
�вW�p���#�G,>I��Q�#!͈�أ��Usc����ۢ�D]�[}̭8c;��\�X�g�T<tk$��ɍ��!'�u�BW�{aEP�g�m�<%�O^}�$Իc%�r��XU�?�b���Y\�F��	�R�Z���� )L�NJC�՝���U�ݰ�d���:HG)�G6H�o�q됹���Xyh��ǈކ|�L��~�)�0^�Aж(������[�D��a
�Za��j$��T�_��o��ٴĮ���U�H���#W�W��.���N5�D���Jpl���k�6�}B<�2�W��s|a�B���a,�īHp�}��6�gg�'h����A���7΄C<A� $�hkk%�7�4![�w�������Xg����z����wa�P a�b��#[�d�r���y��`����m���"�ejY0���JYF��4ƛ�2T�)�(\��-�.��ۖ~Y��$>�m� �5OtWu�aj$<"_�AC~Gp�o[����d:�����:o�{��o�T%.����:!����j���E�a`��N�!��3��;͈11K9f���_y��}z�@�"��@����I�_���kBȔ%�����L����L(9���<gf�82�,g7U��S�%��tIC\|+�E��Ց��X�d�1�mm�{�M�"Y��Y/�!i��{{�,=�J���N�?��=�҃�$������>���_
��Y��=e�fi�=pU`r0X��M���m,�$�祿>��N3�٥�Ohe/�ѕ�,pt_�~XH�~���bajtyD�vmv��ń�䘮��ǴX��g�r��a��p����!/_K߁�r�V�W�[,��ߗ�}wd��E\ǯ�(ɷ}lF�xg���K2�@�6�r���s���*�c4��,y|��+O��_L]0�
��f'��.%���2�O���wխ �\�É�A)�[�,"Ƅ�����P��A�e!�� �_g|	]Q;(IM�dжbY���)����W?U�-���E��[P��X�Bgp�Z����ߘ;�l�bX��)D��%(�޴��{��۵U��s4�������@�vn�]��;P,�Ki�a� �W� z����|0��΁���o��b�'i�t�@F�����2��������ʡ�FjR�'�'��@�܂�Z��f��n�����?v��vm�T�z�7W�6�0U#h���]��Ũ�`�]�؊���'ܠr�%�!�)���\��P�.y��+�x�+Pw蚛�r8׀n�$�ףZ(�N7;�U�0ɜIԙ����J�TBt}��uw��Ѽ{{4-�~'B�o!�^����}���2�� �GP-����PI�ر��/=0a�[�� J��	�k!��R�U�����������X��ӕ�	�T����Il��������XEp�k�z�vz׭������Z4����]ɛh�Q��e���c�2t�ؿ��
�g�l��=G�U.���W�w��ڔ��f�XO�պ^��T��TW���!�w��L���n��J��+̾� �P�"?ƹh�Үz(�ۭ���m���]��(]��H�]�����ʿg<�#^�����Ƃ[��:�TYC��֣��:�۝��-n����3�CQ;��Uo�;��	+�ר��x�S"QSJ��|6�v�h�?��XѰ�?Q�,5��iA�,n���p�f�?��Ӌ��[�d�G(0qB�������)D{3qB��Cv��~%P��g3�C箄h)�z/X��%���E]9����F�Z7�O�͊茥�C)���L�$y|Ǐ���'u��O�`o3�>�?�&�����۳Ҁ_mvoD.�
R c��\�8�_��Vk%��˜a��g���~\ON��^`�����r6k�N�hl%0�q�$Q�S�����Rך�t0�0�Lɲq��D������ ���P������tՕI3�f���-	��d7��@tf����R?fz�܆��H�u����xt����Z�7c�V���E�}uf����fR���?+��9�(,v�W� PD}���z̝.���k|� |�"��4���1OL+S2��q~�>F&�����s�o���CR�#��:��d���C&`4@YWgo�jx��>�a+��`@u��勫I�u=� �!��k+w��-YBb���И�&�*�p���Y����_ړI�N)O��R&��U��X^��T����q����>����٤�;�ъʊSt����'(�łR�fL�R�3�D���u��4�A�%�Y�'a�~2��aepx8/����AS>����/�뜿Yw�Ve�KdϺ/���!�_�`?��Ʌي��V2�`�P�t��G�<�D�5�m�]?���Ϝ��B;���W�dR�Ｊ��FP��?w�㪽充������u��l#5���z}O0�L�Yl��<ڼ�����֚�G�(@*ħ�#��S9O��m��P�i<��e�5e�ZsR^�@�]��	��C�;����tm�!�2�1���=��1 �R�l�?^�d�^I��0���{��0���751���	E9��j���^����G�ͳ��#�K�:�����Q�Rxo���6�`Q��7���j)ѓQ�km�\�_P���;|B)������
1�����8��'��$͘�;����_.��(�&���籭lU��A��x��?-��d���8f��{Ǜ{l#�W KǤ���d=�hYlF\G�]���-��$.'<�qyZ��#���cK����n�e�VvU��	�a�W���'���|�@z�[C4p�>��n����x�!�I��X;6ٛ*Nc]C&ʘ	�Ǩjr9���ޖ�t�{Ϊ����A�ҩܮ���WgUj^��e�����¿b���:�	*��Y�r��	6��g}����2�l]��&�;�;ʱ�~*��K�3��7Bct�/��:�n6���3��%��dh��NG�y�#�2�{�v��>��VƎP��a/<�&��� "����
����ER��\=Z�l��l���9DFp�!�·�%���t�Hh[@5�Pam�vT7�O�7e���hR���rܴ�OCZ�!j�i�`�"=��j�*�!n[ؐp�)��[S(C2W k腘��9e�<����޶�$&O[F�4�Wы �ϲ&Y�\g+C?����_r?nRU�])|�?��p����H��9'��Nմ@����]CE���sK_���1�D@`�$��=c����T��dO2/���.�X���[����Y��S�8�Be|�jY���c�^��s�e8�r���5w�&�o�Ⱥx�^�D�,��s� �h҅O����_&{D��*w�����0 �TV�!öD�"�y�psa��2(��Jf�fi����lh����N�٨b�>k١^`	d�1 e�[�*P�� ,W<q��Ze�q~Jڑa2��w�,�)��*H��l>�G�^L9T�Է�qh��k�Ɯ�hx����O�N3���Le������B����4J�T������\F�*�lR���m����jx�.��V��ۉ�,��EY�;��k�9vN�V�k�X����R���p���WP�>DYGړ�,i]W��L�Ɲ���lߒ�����$�>���ZC+o��gi�TC��(�ÚI�����>�{5+��8&YV��U���`��(��� ������s� ���C��an���mj��-�h�`^���������<H< �ut�0�ժE(Dq'0R���5x��Ld+=7�%�s�=w,;�p(&}6ǡ)�
�Rkv�,�E!Ѵ&�b�N�ʾ�]���<�R��PO��k���NP8�˷����]�pw�+�2?є�8H>�f�H۪TB"�Aȳ�-�ʮ4s*�&#�)�Ԑm	r��u'BR�J�	����^w'���"��	��<���p��i䁒��1�?��'�P-m��3ʮ�0&�8A�"�/ ���n��k��Y�O���o���G�zr�gb�
��21����&_\�c&!+I�2���5�I��H��|��d5�:h���$
.wE]2�%	Սy��*��L���as��u��d?��b{e���s �ѧ�X���#��˖W^-}�l]�$����<��F�D�u��΍���}Nw��˓{s�Z�#�hqf{�gf�"��s��pY��ӯ�a$�C�kkuMVչ���E�@L�h�aiI��]/��n?+�-��;G��,�Ƹ��x8�HӹeL����US?��P�2CS��7J0��NS��슔��Cy��z��O)u�^Y���q�%��7B/]@�r���Y�h���񲟗=�ǟ���ɸɜs>�[逴�qS|U9���g��W^�M��6��}#��0;�e��|� ��t��,?�W�zJ�{n�鐷;}6�#�h��_��d��&|�ҝ�R���5Ru�4��(���!k �]B����W�=�ƦP-���)p�������3G��0Y��`;CV�P �~��3�f�$R���Sβ����.C$s���IVֈ8���O S���ǡ8��LZ8�b�;uFfG���}d�sV�\܀3[/V��$��帽ZEK׎Ŭb�`�&i�zt�%�uRl�|]��8��	3 �<W��l�DW����`;`2T�ڟ�����Z��酊E%a� z�Iϙ��d����P�kb��,�b�2I��Q�©�8��T3/�2r�8^2KVY��r&�є?����i6�g�x����x�8N�YnBȮ�߃�Q��9䉻=�6b�&Υ�Mg����].z ��-�Z5-����-�L�ߠ�������%��h��yͣ�k����K;�!lH�gb\�b��ƈ�AysH��.�RFe�jr���`�F��@шb}am�/���V���{����z��Z}*���w?��C�"�k%"&cLQ_	C�0Rs;�x�2!Ϙa7!6���!�)w"����/ ��0ԴdF\���E0㛦֔�*E�Uw@
�3X�YK�&�D��fBlq�(L8I��ih@#'~�.�H|	�)��QMH�%Dl���[3��|�!&
"�iU�eYH9q�$1	�ᆶ}�PeV�Im`��"��Ė7��񪻪��N������<W⣚5;<G�_���ԫ���$'G.�am}�>n����j��2-��T�Q�r<��,��E��Ѱ a.6��#���qm<�<_;W��p��4e&iq6�����#j�їt`y��M�@X���B�K���`���*�����H�Ϻ7�D$�K�*�i���(LR��S�AW ��zi-���{XgkD�i�^V�2���=�pEva�Zj�#�m�m�`o�V��T�t���r��i����&�1�1!�rľi^�6]�\�m[����[��Bd�ڝ��v�۸�e��J��l�b�e�L�����z;�z�By���t`�D�T9&Պ�Yop�������TS�qy����b#�8[�k����6��/x�R���8)[0O���I��n���m����i+��u��dp����J=�C��L~#2�c�Vyrow�5ح�.���8����6�����?�
������B���</����;�4/�$S����-�� n���1�L�۳^��W�'�'�Ml͡o�2���j�u���t�P��3�@k|�t~���1�|��DE�R��H�k�)N;�s ���E�-/	�O�l�o��L�����:�	R�ڲ���2I�s�"c��q�K�G~*k	x���?��ԡ�?�e���z7��e��6#���BE�W�Q�vF�}���/
�%�	�Z���},^���]��5A�ڠ�qUз�^�i��������_8��O��J]��aR�Z��T��eԤ�2��aHa�]�p�#2��M�\�����<��/eq_�EB���]�G�Ⱥco]�������c׻8?��鿬��bx��� R�M?P��}+�D]ш�c{��"�5Ɉ�]_��{���MW#V2����~��bgPV��a��NP��)��*kĂc�E��0�iH�K4��r�ԝM^Z����n��]ăv�@-������|eJa�'���Ё�$�Pg������o2������t@�O(�|��%��H��p����m����b/��w����;�W����ݕk�ޗ*U�)E�9�g��G�J���}�pF?�@�^;�ĻWCJP�E7`�9�>��j&oawG����ʇb�7� c9P���d@�as�t�vCJ;N���|���gS��	Tǝ��v��+5�g�N�v�������3�W��Z�g��*��r�jc.*h�b���/�+{Qǃ�U�M���r�c�V�gm��v�=vu��>�q3!�K ��}}�@4:�M�¡"ۮ�SIO�w�&�e,��^���Sb�S��cC��tHQ�H�Q�n��ܪ���h�v�7����!�3Uc�GL�+��G-/5�x}�!��ꊒ�x���s � �����f��N��E�]���X-���h�5�\z��Ng����`�������_�6����\�����ͺظ���%�<�݌�7��lQ��ֵ��Z'���pE����s��v� ]�OmʶJ��u[���
�h�̠����=�f*Q�CV|zg8Q��#���c��A��G� �ֈ��TY��� ����6�O�C6;�Y�,��ѢRI�0dE�C#u>��ץ��E`���z�B��|R�tǌI�4h1�ܗи�瘐3�L5F)����&�w� !��bl֒	��$�3��ϛT�\�
e��{z;�6�*��w�uM�y��.��� e�&5T��vT��nQ�Á� b'���B"(��Z����]-ĤįdkᓣYՅ4)���N����P�ٸ���<�ew�[	����z�V� �f���Fꙣ���r������/����%�,UCk�lb�y���pYRUE+�O���*�� ����]>9�׫���j�����Qm����^��t0�AP@� ���Ҏ�&�)���f�/�՝ֳݦ��1U�f�|,��Y����>�U�Z��E���j���'1i�@
}���n��x��[�����ͱ��^x�3�~�U{"V �n�*��������}�n�1v��.��i�I��@:���* ᾨ���vT}�j��.������.����'��T�L>�?b����Xt�byMF���r�����f�UX΢�p�T��}�ޭ���2��MV�D�������MJ���� 00	��HARU���]��e?���G��8c��l�������ެ7�es����bp�%�C�a��s�7H�-����S-��?~Q�J6���U/J}AEh�7�}:躨w�yQ�xy@(u��=s�ng[mo��&������E���rv|�W���#d�l��F���ݴ������(�4�y��߷���ϓWJ�5в�˰�Pv��\r���$�Ԓ�O�xO�~;'Z0]��CD���LM
����3<D�~aD/�o�m����;��Nr��h*S'���
N�e���e7����h�����_�Ac�gd����y�ǻC��F_T�[f��_@��t�W����������e;�QZ������`�{�ƣ�N�9.ч��b��=" �i�N�O�
���;���/O%+�}A�����Z���C?�S� rQ#4�/�e��8��WV��`��>Y� �3��4�`�v�������\��p'�	�k�ٴN/�/��i�CpT4�������<���z�;E�Y����s4��}S�İK]�*%\=K��*-��S��u K:�%�Ȃ#�g{@(�L a��} k�nD��sާ��=y9�k��H�*���`C>�=Kh��S
�.]ږ@S����N���R"j�ڳ�s��K3��QD�ژ��dJ"a��i9]�4f������`p�E(����g��X���A������L̕���T�m�����W���D��EE��!�~���*w��xu���O*t��+Ϛ�+���;1�v��6��SxsI]7/+��	�5?M��a�4��Zh]�,�cOc� 8��_U�[�MCtgSRq+�w�:�?�+�
���fϘ�x�䪮���	(b��!Z�[1��򺆢�6��Y�ْP�ݓM:���\�u3c�g�NO�F����֮�F/�c�v_J��X8V݋��-��������r7�Stw��ڡ�bk!%ܨ��,����6���[s&����Ah3^cв��E0�B2٘]	��W��Qޜ��`>�3��V];�f:A+S�%\D��p�)�aoE��DQ���3�f��1W�g�D�����<�=@�/�h5�E�����+U�JH����
d=�5cȚ����B�|r
��2N����SF�437~���B�!j�m���_�*�Ҙ��p��!If�¿|���H#�&���l�c~b3J�P��VOv�����u���FV�6o��'��D���]�g&9;�L�j��)
��f<�Ԃ'R��\���Rc�E ��	c��U���sq	��&c�u���\��m4�nz��x��#W��+m6�}f��>ձDr�{�ʉ(_�2G����nZ�������?��s��\+�P���0�$4� �����g$������!F�V����ܲOVӪ���:���-����X�ތN�y .̈�C�Ui�|0.9SȹFR�\���$�WZSѨ1�UP�w0*�Fe�u�S�d�d�����M�X�v�C&D�>�aN��{LK�+�[�&�$�u��B(���&+�����˺+���%�˃�i;$�."��hI��4t�
$�A=#1�vTp~`�!�d�SG�$bYQa����F�\k=Lx�����]��E��c�16�La_��X�g��o2V~����\d����!hCĸ8([���j���ts�8섘]�e�q����
�>䖓�u�<�Gev�'g!7�=�����|� �⫘j
���^��9�$��u��f8�wm0�k�=�dJM��!�a/���Ja�
q�?������5��n:�I�#����-�LY�6Zg��oɤ���u���M�A7Ec����`�#�N�����(w�鑠�b5q�ӢٌQEu�C5�UМ�M�>�rS?8���8��B��O�� b���o?w��k.��F���b�#�s��Ȫ�/���m�TFU0�)7;V~���m��>��ۊ5�5�X�,��t��ٍt�����v�� �vg���&<�TT͂��݀R���
;CV�f�L^�ތ���������U��7BU���x�R���Q��e�Q���.3��0���QT7��/3-bM6�t�
�E���/yQ�y���F_!��x&�͙͘�>AY'�Rۼg9�P�:��F��ټ=R��QT#��}�֊�67���Cw�e"	�׭�l�}ˮ�f�U�Nr���'�KǗ���j ��t��Nru���^y�)��[Y�쏋#��7cϙ�#n 䵊�/�dj���o��,p�U�>�։{!1皮%h'�]����*C�_���"���:�O��,�my���OI��F��ʝ�`OiQ�Y�����Z&%����>"�fsh?�h�D)�$C�d�)����Ilf1&܁�o틻���d�-c2�6�=��韝��8=a6titI������`+\p�x�S���e%���a��.�`�h�r���5�>��l��K��� 9�-ǅk��m?�Ϧ�9����{bo��ǨEV�ci��ˁȥR%�ebQ�$����*��uJ�f�Tl�_B��OH�ԓ�ޔ�&i{�����ݶ��uI"�5�4�7؆
U����A���&���2:e��}����9��)>I�N�7�zP	�-�˥$��E�+��.�WU�N��b�J���X0�e)�d�%Z��(��������Q�DK�LCO*�z�?	�cNG� B�Z͈x,lCި8�q���ws�x1��
�9��,6���g.�ԇئ�BpC�GȔĆI>�v�aƵ�����o��q&���Y?�e/���'W�c�3�X,.4�r�%K��\�A8��$���2��$����&%%��Qb��dD3��c�M1ொ��0�X����lݎ���H�w�V
18�%"<�8�(UZJu&��+�Y��P�����I�<��4�F�������.=�3�:��y3�g�p�F��9I ڦ+�N��n���=J�������oS��k�λz�|K�|��`�	Q3%���Ms�(�[����P����B�pЌl�z��ING�ܝz�^_��.��!#��D�Bp�x�fR��;So#[�,��3^v?8Laz�<�G�Ǫ����o~׌��_f��>l��n�3�OV(vmԩA��Ms	t��8���5hІ)��c~��LZ:���m��#R8�������53�V�y*RתQWfL��͜:��TJ%?���� %�td����upG���S�Mqtx�@�;�mE���w^7\6��t�v���C�%r4��Á��+��PEC�8�Zxi��sܗ��qs�h���Q�j0=A�x��ψ�-��l]#�Ƥ���8J������� �b�;�;6�P�TE�8�}�;ӯB�(���[I���!������I��mղ�*ժ7����g�Nn�]E��ܭ8��	p?�����E#_�o���6�n���`+��}E`Xڅ³�G���Գ�#�v>c�;�,|�9��n�,N ��Y��'Ǣ��Rw(�����P�X�s鴳�@��u)��U�~�-����oG���]=��G¹'��fuK��� �vzj>�p�X�e~����P0p[vX(��6�m���}�Z4�b~i/N7�<d��_���_�6���BH]+�AS���b��R%I��mZ�;���ZO�>��0y�v0��W*��������3��7����	�?��ͷ�R6��_�?����G�ň�}��'Bvn5S�q_��t�)����c9Z1����T�G�	D�Sx��Uȉ��Z:&�����	є�2ɹ���b�YR��:���j�p�݀~��㯉^���C��'�D��V3t�Ѽk�2]C�À7LB�ߦ�e�$I��`�sD尼�0�h�Z��9��jG��־���ѳ�x|
 ��A�yV�3G^0�k6r�	�^����3}_C�\o`�Ի���D&x�T��r:�F�?��LmXt$�vY���	�! �)V e;rp?:�.<���<���2-
�Z����7��f�򆼝 ���Gqe���q���U{n�iR�ItW����O^�1�>��yW�=���(�N���6:�H�e�P�=o$I������F�~P�������/}>��" 3��+P�˚��/����0���ą�t>n���C}���-��п&ރ��k��Ȏ7����P�f�Bp��տ#�CAFʥS�߽��,�3g����UJo��E�:��~��'��f�RD���N�t���@-�����}8C-��.V}���и��ER�-�Q��A�N��n�0�_������`���yu7����SP��bUrEb.�[ݢ�յ��T��7r>{��`d�K*3�R}��k���w�)�LӉ�_��%��~y_��s<��!a�{�Y�����d^܈D�_Z�
=�a����E���h�C��,�Ĝ��*P9�U+���J("�Q#HW��q��FK�4	�)⛐��F|��pP+;�]|��9t8��()�^?�u*0�7��PAy�{3]�f	��]~�-K|q�D�|���cĮ��L��#�9�:��Gs`/��/���{���1�L<A���N�ɂ�Lt{�pnu�1=�2�2��RL�H10��r� ~Ex���]���#�^�����L�3�2��G��H%|L�#�pc���*>WQ%=_+�����;��la_ŉ{,�6���(�~g�?��N���yH����*�@���1N1�?+"wΔ�8����NO�߀o�e�"FS,���?Um�1N�^����0`樝�fV�h��/���Q����|�k���N����[������Ѵ�I]��w��X�(�;o�C�n&Y�� ���^��w�ǽ�.ӝ��6@J><��)�g�3ah��|���E0{�ư�b.������s�Ho�E ����N����hơ��Bo��l�]����ͨ��W^�{��쳬�oAC��kk�D���l�>�̇�yOoO13�j���?�"�b8����xJ%Hc�����bv� ��y�,qǞ�����/�Q`B��η�z�}�v��D�#�q�T�f#�bcίS=�:�����Ӎmr��.(�*_S�M��<��r7�V��7b��f�8R b�M��l�c�|xjνw���V�f��B55G��#���e���m�\����s��c����.���aŊ�9E��$��-,���>t���_ؘyρ,�f�\7_�����K��J�|h9`����ګTu�Zf�D"6����A�y\vV =R�[���%m<�`C}oYĐL�Fb ӔZo����	�L(:��_�����9l�(���H�j�����'���灧��zP��-e�&$r���q�T�� }��N��G�Ѿ�U����n�)��M{��kZ���a;�:������`�a����6�Ejm��B���������VDk���=��'K�����+��\�d�m�x��5���ൊ������ ��}Y�����.
���j�+�f��KWa���
݊����s'��j&'~��E@^�sQ ���kCH4�RHfCu�p����?7F
x��[V[Y�22���UgҐ-ȥ�FP`88�3�M�D��LO5&�P҆��IEJM�Su%��Z�+>@�# [������6P�B}؛:�G��'�z���Gǰ�����-�/]K����9v4T����LJ�+�?�*l�{�΃�E���
���mM*^����_���Z%)����t=�Io_L�v�2������̈�G\ܯ�5v��4{H���q���p�1[/W�_3z�/MX��}]�����9��y��6�Ne�$��JF�Qj(jd_���8;>$�}���`�ݮmL�]��a�.辔�����;�*��~d �t��]�~�9x�����V '?CY��~Y`Uo��c¤�����HL���%�M����Ǭ0^�1�	H �܋�E1�O��
���Q��Є7\���)u��w=��jlӦ������#��Z����3�П��DzU���^������$q3_퐏�&��λ�B�n�%&�m`���mum8}����m*���z���mYD�Ř��bB��t��~u�������l��"<3;�B]�]q�/�o�\|�L	��)pq$nOs���K�n����������pl��]�������E����9�,ʹ�=�a<ǀ���sR �&������y�,D٥W��K��\	:��Ǻ<��W�v@<OĎ�ԡiu��`�j?�u|u/
ޤ�j*buí���.�84��b#��F$��>[գa	 ��{+�膧	��O	�>��0�����D��5���X�Nua����)�]Z\���P0��Ԯ���!���
,�RZ�)>�*|*حcL����eo���mM��!���<����=:� 0��3[�P�0}��=���X�6oF5l�Q����۫~�Ei�'���u�T��KŬ@�3#�M|�S���}�9����!G�R(Ǆ���\x0��HD�ײ��W�D�B��u�a�ׄ ���Jpj@�G�C���ӓK�! "Bi�%5�O�9����j�XHϛԁ'K�j=���١��<��ໆ7�mPX�>˭V�{��R(�k)8�)�|�-��/��s[ݺe�sT�^�[��i�[���~w�"�;'��|ydg���:�he��`%��ւ'�S�c���>h�x����vl��ۣ�2�Dд���{���s���P��*o�	m2����(�t����J����,��p�w�le�qT�tz���+�T4�H��;��S��\�܆|� �n�]�����9/ 3���f�FX'"��[�x��5��I(��\:٭�Thd��fbV��	��O,q��u��X4W6Y�)IW���ƥ���#l�� �U���C?� ��X:MQLQ�� ��Y>S�@>زG#�k�I�F/������������I!�A�E����5�IAX�����Q& �R���]Yd�Qo�0�U�զ/�/||5��*�N��׷�c��Qڥ�D��XU�d�Q�L;���gם�Z��qvY����q�ʖ8B�ɳ�c���9zӨ}�8^g;.nE����A��k׫'��ۙ��S>�#Q�>8��Y���RL�TFь+S�H]�)�p�nSF���uZ1'tџdJ��Y�P��0�j5a��`T�� ��
��ӕ_�1�b��D��t������q"m����|z�s���M;b�#%m��Pܺ�EyE��|D|���Ay*b��u�Z��*/�aL����o<�Vx���)@��G��OI����젟�p����r�Ú}������0��ے:-i����]�U������?( `��*���c��h]A�����f�����Ds��E�������z�
JY�3%�M(��\�-B}���](㗂��851SB�������(�X����\N'���=�i,�5��sv%�LF��hxM�̏�� 	�p>�n���N�R���B}7�ujb�	G��IF�����|t$���6�΄s�H�I��4�20�d��^�����0�p�E^��+8�1��&`��ȩ����4,Q^k���p>o
�r"eX�C�-<�	��Xǥ��. ��P�b>G}�T�I]
O�\w�h�"qP�f!�OeKx�R�^b,5/h�e��ʾ�bD��䵃_��c&��cآ��L�~��X�9��2�d�Rs��e��>�3����bD���?f�n�O,��0b��h�(z��;�թ/;�L@��&e]U�7%�A:Z��ￆ�ڃ���mݼ*"i5����'���E�P\lP�흳i�uf�>��z ��:��W��Y\�OJ}��x;�����9a�Ey��;�ԯl2	P��� �.)�Ge@��Q;x��ދ9�r��mN���S[ylv�^��r�C���Y��翞c��Q]��	��t���8q��3�w���x���$�+��7�"i��T���f���<��I��֗a��D۳T'�(�WedFJ��2p� �I}���h@
�T�UC�
ONE�qUa%70f���L�st]Ë���7��\z�q%�}c5\r��+OŅ��XuM�*��\K*V��ָ��-vM@��WO�D��*
����*���*{y�~�J�A��|/��X��%j�����*�_>���BR[d��'�a|�j�|(}��,&
�e����uVN��9��H�.�ī(��Њ��B��ƿW�j[����3M8�`u�H�1��'ț&����LՅ�6�I�D�lY����m�H�.�9�7rJ��Y�O��m�.�Ŋ��l'վ����yM�IQ{A9a2�B�ڀ^��1���"��"�Rè������w��FBu3�$��묋��eeȮЅ�2���l�������q.Ѐ�t]�#�4�A;�� ��-!����v���y��F6������M�ԑ�����Y�8�_y;~���q�F�����H��k��NJB�Z��eo0�|�mB��ӑ��u�n��#>圵iИ��S����4��Q�voJ��~��d�T'�f	�,�P��#�K�;����%Ùӂ���k@���|/�R2��i[+��C;A�'r��L���4��,���pOz)5��/_�o�_����	G�E���OYhE'����%�/H����p���R95��7>j;	@Q� ��#�IɆ6��hŭ]���x�492��&P�pϢ�;A���N�	,���3A�d�on~7oj/�R	�#b%wHSF��2������!�����[�y��
1�@�s������<�� T�JF�{3�(0��� |9�fM���1^S�Xe�7��	�c�7^WK
�>�l�K2TA����M��Z�%9оb�%䅛�a\�eq�����6A7Fwl�>����=��KU�|�f���a'"kՁw᎟�]�08Q�mw��\'���g��ɸ��+!��	���]�E՗?p��u�����
J��<�'���N]T�X�[�DL9yQ�3�vD} ��s}��P���I��p,����Ŝ};�t�ǎLqO���nr��-7����(Ci�	Ƶ	d�d[��[��5��-��[�>B�+R�Wo�Bܦ%�Y�.��a�o�I):�B�����J:��a�V*zl��� ��\�p����ge�{{<u�Q߁��o�6��4���f��rʄ�z��,��J��k�B�#�%"\(�`X�[�}5b:E;,X��Y;q�A�{7��g�~2�v���T(W`��_{l��%��D7
�}�}���3a~�C��'J�� {z��B��R��g����E�)���}��>����1����=f:�d��H�O`@���nج��#�#i�&��������p�6��Z��mȞ�=�{��d`M��r�m:��C=V�u!k��T|���H-�woC�7x�e������� ��M۝"3��6���%.aMUh�N�De��j6Pό
�|�{�	ޓ7��LX���N��:ݐ�=Bj>38�Xܘ�R������]R�����ݙ_7P<"�>�)��O|ӽ�7�Z�a���Kf�GM���!��L��UeC%���������1�X5y�}%�X$ql�s���,�]j���?�(�S<+�k>��� ���A�x�K%_4�ü�8�	�MνC�1}	��<K��^3�!�F��3�4�G����j�Wy+o�#���?!ݬb|>6�hj�ؚ���N�J&˗x���Z:�A*<@(7=�c��M�m��0�TD	���s-b� p_2V�������Їo;���yj�����sݵP�po�o�,�����䡈f���#���=g/z�;������y������n��z{��T�<lRv�d��+��;�]��	�I����ЀŅ���sN�Gp�u��e�; ���~R����D���u�@ {Z�V�+3��-e/�`g��誼{�hS6�ǭY1����A�Mj'f���8������Y»KN�z�E0�;)�c2Rg{a��S9��	�����!�P8nj�T��vp`�P��K~u����_8����)lr-廭^�S|&ں�H˸�Y5L�#�����MVˋuN%���}=a�Gl�mxc�,85Da����C�`	o���������J4���>и楿 ��+�_��t�zN��;m�۽ʽ�ƴ�(��voh�uw���7�[8I���|7?�m����ͼM���e��.���G9��Wi��k��9^3xQ�$q;?�+O08FG���<����R#0�	K�'O�8g\����˃���n����*擼�0����Ke&)lӟ�֯t0���3�|�;؝�Y�#�Ky%ǧKC��y���M�&A]ʾ��a�Js�x�R�b����T��P8�*��"+�X�_P�LdgEO��!"b-�&Z�D�^Jxv%9���xG��*|o�/��<ыB�:� �҆�����
�y�n��e"Q��li���x�@����H�~\���$���Hu�C�!�E�;8�b�����:hI�5)P_0������46#��~�C�H����\�0�>)4p��S��Z�|���{�'������|�VU�����rWW��މ�(��맅H��l~�p�D%[��{��2Sl�u	
�8*��.Vv��/jB����a��D\�U����q
��B�ȭϑ����ט�l�:Cl�b�G-�l��npp�4�W����|��l\F��=|���	�=��Vs���E��d9 �3�jzT���i�"4!5���˥��,������
cО�:��<v��YGt�i}���^��֥�鼛X3���3����Sl���rK\�/���g�Aʹ�]~D�}~�d52;g��;o6�B��7�~�MZ�
��i'��p<9#uo�b4�U�)�7p�aY��si�F���^��B|��L�>>9��DF)@�8�>Dl��E0P֡�*`�[�����K��?OG��@�qh����od����>œOv���:{�-��6j��s��}�����)�3\�6��Gǐ����澨'�f�ᢀ��^�xh"�x��y��BǉǱ���griC�js�7\�g�
H��PCÄ��֙���{
9n������%����Z3�W��n꧶�����1V>M��Kx��
Z���;pӃ&?.ag�)%J�#}�HE�	ਠe���o7�&����j����z9��h�^%?�>ݸF�7 ����0O��ݜ9)L젤9��a�4���e/q��yɓ$L�&�bt����]T��վ�#ǹ�<���xmk��!�fK�(��fn�H��:C��q(�R�ȿA�Z3��E�����5������$hž_�A	��Gc^��乛�{�o#�DB(rs�w"�%��_�} �� s~�z�����Δ没��%W :"3� -�1��A��gv��"�ѕP����*҇��G���§0O��3X�e�S������P�5	't3��K8j��!۽F�����:�R"5�[JN_�΃����!�5��'�?�L:EPB�^6�'��OA�s ��.~��z*:�ɓ�s�b�a�vPOv�\�G֛�W�p��(�te��;�
o��z��6k��D!(\p�*���F�X��=C��j�NB�n��w����Q	�������S52"|�ny���hd�����b���&qJ@/�)���:�HtƏT�`��g5�<f�' �s���~|>�buް�*}�|����֨���Z�ɏ���W#����%L��EYùy�2<ŪԨV���������Q��|���h�FF��*춥�G����Cm����ž�ɖ��,� ��g�ߩe�+
$����w{S�cѦM���N1�[#�ݏ�j��a��C��`�wfc ipz@CHQ��!���/�1�W���xk�h�I����������`z�;�?_7�������bJE-j6(.y�K�(1*��ˎ���q�T���f��a
ҬcV�J5n3Ƥ���ʪ u���uـ�+�|�$�f�p��Ou1O
�gߔM �ڲy˭6&t�_C=�>��J�C��s� 33��&�9RL$�H�,��u��L��g����n��$[�B�!��S#U'�5k���"�`l�F��"�*ѣ,cS�+35��uC�Ө���le�=B�a�ܭ����Y�_9�����.�#��8��qZP�oz�&����?L���"?�GH��1��BR?�c�#;�;a�p�A�*�Q��p�ڤdK�|��铪8N]��5�.~h���-qC���z����g6��su�x��p���+7��Z[����%�ɶ�#��g���ؐ��g�m�n�N#/۪[�y��G�Jq�����jC�g�baԗJM�:��=x�C�H�9 O�_f`�W��<)Q�S��3X%lc(q�^l?Ԡ
UEw�����,CX��b�sv�S��B��ub�p�G{��a���4�>,zgG�{(FJ#�3��:!!�U0�F�P���M,���(&��]<�х@���MM7�����?�X"��Gk_R��1��;E�T)��`�Y��z����7�сH�0�W�|�f��T�g���b�M�
64��V��F����oF�z8����a.��G"�Әe7/���Q�8�y�C��!y��vU;�����>�3w0 ��u�����Q�z� ��A�}p��jpOD��0�z<Ф4�XZ��o�?�$\���ɶ�p�����"�������$�X��ʉw|O�@e��Êto����eI^��e�ƽ�v����^�nr��~1m3=�f-�����+�6�\u��	7�I���[��>��C�����>�����&7������:Z�ھ����ENY �AQl,���Y�b�a�Q2BW����6!;�,5�3����?��&���[Qvld��9爞����\��?��rd��D����Q���G�%LM����ɍ�Tb}�$i[�g�'D���85DSQ�_�� m�2�{��b
��M�\1UX�~������Q�R2g�"�^��`F	�m���9Är@X�s4�[dDt!�#�����B�n47�#��aW�\%�~��F"�3Ʊ�)f��[	L0�<��^{�4�w5gq�x"��Rђ�:Q� ve���	Am�g�z�|��UӚ�s�R��-�|�Tx��[v7�����0�S�ȁ�O,>U�����Wy������_V�6y���6axӱV���k>�=�M�/�����e�%P}2�0��,�.8�1�������xi�t�п���QB�����ְF#}��?��B�S��>�2٧O����G��BB��t�pc�G�4�b��9�bq��{9pő����"�q.9[w�RΤ�ݕi<b��*�@���G�N� �"��=�+C�6Qp����6	�-�c�e��3��ˌ
˹����p���[�`�F3�B��:�R�g� �޻(�{b����w��r���uE��Ɉȃ��	�w��|�]�.?ޥ��:bWK1vK���ƷEs�?8}b�������oG���NnfksE����	�&h.i���'��n:{����{y�
�U��F0��UFg$Xf�&� 'T��Ga�,�+��T���*oG��	��9�ֱ�l1
�<��eCȻ
�a���y��)au���Z_7.ɒ7{�c�U�
%��-��\���0'���$�l~��"I��)�Bl�I�R=�,��죪)>�vE�ҙ6��X�e�����`cV�z�6��Qm�����@���o����6J��%�Sg������%c0,(oȊ	p.�$�B۾ʼE��������Da���0�6B����Ol��� h�۾E���]w����@$��sqA��I��y,���w�̧YDKQ\�`�������>:������g<��l)����Ue��F?RBv�q��@��3�<����2W��K~�Bb&K��<�l$� ����J��iQ��!ǌ��hBɔ�G��¨�o�z\b�k�Խ�@�� n<�w���w�0���Pʳz�>���+�T���>��HVm�nsΉuN�'�Ǚ�#=�����(�!�&�[{h�"�Y�����!��E�< G�ɫ
�1�F��"���><��lz8�/�1����t�L�x;y���4�o�G��H���o�X+��qD������
������n	�c�4�#�*��L�ؾ|Lkn�c��=���4��H`|?����ߚ�~V���+5�y�����k���,,�}��:���$x��՗
;Q�!���x�M�v���^9�X�A*�^�0�N����oj	8��MO�F3m�>R����E��K�Ԍ�͒9��x��s���[ a�ΐ��5�W�
ס?s�+��E���nn��d� I����:�I��F��kj���(�R�H���!:1�v�����$��`�=+q��ͤ��e�a9�[���I�A}\�%+��l��U}�u�M
qxd�`�0zd�i��@�m ��I�]�֡�"���R�1ᇡ\t�L��k48C��F�x��6YF�����2�;Ch3�l�����[��j�/�<fd����������1���ң���f'�[��1���ϲ=���߹��phX�������E&9�?L�i��`_h<���<r	��ǰj���E�G:�(��8���޺��mP��J����"kP#���vpb�3��`|���Z��,�C�g�����U��0O��Nw�3bkV�S�{W�0�ؕ��7�^�	�UZ��E�C�&�0p�����F�u�DrlÂ0�����dr&��J~J"��3�׶���+�x���U풻+�^�|X�.zl"^�E��'���͚�8�
teȭ�&x"wڹؘGr=Ė�����D>��Wۂi��l~���ٳ��2����,��r���k���g{s�$�ol;�qX�;.1�-�'M�z� ә���Y�V��-Nՙ�a(�'vĖ�>Ɨ_�|�%Δ(�V�(�x�v�����Dׂ�D,���05�,�;說�S\���i�p��l|�x�h4���G��a'�Ukw�\�&�K��R�]�hm��Vn�9�\G�"�Q;�x��i1~��q��Ho��z"�?��G)���5}�`v9�0A��vot~���hǧ�W����:��	�fo���v��%�0��~�%�9��{���@Lz�*_������h�t�	I�V���!�SߦK�V���=;�H��|�u��������x��-��G[7g�'0`�re��^�X�z��LmB��Cp�{rsm�K���U.śf �XL�o� 쬱���a4t��a��!*w�n"�;y�,�k��)8(֘��ߦ����n��[������� `TY���5) hC� #Ld�p��ur�D����("(�PT������ss��N>�̷��V>J\	��5��L!P�ƼĲ�̤�
{�N�����	�6�p������/�#�{I�.}@A��_�pz-�x�L YR�ZR�R�BG}�u����o������]B�Ϊ���EiI���l��{�0:�n0g#��TAM\�D���-�P��`m�~<hCDl)�㶍s1�`������NFV|����)���˱m���/�� 0��ǿc�4A���ߧ��lX����fd�7c����K��ly)����u]�?��"�E���
�<�+���[^��xm��/,��
�{�C'��&K��<�X2�@�)��iճ��4�?}1Q� �{^�KFȫ!�$�XS����jsnqgw{l�5�\�Ek��ц0�:�?�iϾ��&Dh�x�86��� c�\sP~����$�����i����2���|1��3�
h�S��������NU�Ͽ�-+ ��;���O|ǎ������$ʆ#�dy(���G!nC�$��}D�������7��k
�]L5d���R��l&>��㚢�<߃=1��4[&HN)���=r�K�mU�Cad/�x����̞��Fg?=Vf��X�hFZ?��ez��n:���4_i겗²�x;�u �R\��<�F�*�uۮS)$�T��E*�O���Ԓ�f�,B��\,���ƭ�ɸX?���矷3�hO�����u�ݬ�5��<�d�`����"'YG���[AyS\4����f!F���ja/�-�ن~Rh�N7�����N;z��'�F���6����1�@�gZ��
�iștA��J�:%D;=���0r�J���q��+���ː	a�M��6�أ��$�*�d^&��}G�(3�bΫ/B�5X��w�Y{@˧���u7l�JQ��S%8�ř�`vw���c�*������{3�Z�t���	L���MD�z-v|�l��V lP��i�ڦ`�O�0sl;���q���V�V!w�*�T?H��
���'Ơ�6��GpUP�oȮ��2Ά����!�x-��� 
C@���D�̕=ΔTd���T�Y�O�|ß �1��dK�BL�cS���t�P��HD��v"%����vn�29bV�*���+|�\�1��C��
nu�!t��F2��i��yB>������9^tW}���Ix��4ͯ����T�~�%B>t�{7�K�z'��U��;eӦ�H��Ŷ�C:���Dw�K���@hII��a��o�c�����BN)#�B�peY>�DSz�O܊Z�"�ަ�̋_՞���B�z:��c6���د�tʄ�S�ȡ� �j]�;m�x�%��E�	�u,!�v)�KQ��Do��X���Ը����Fc�m�o�G�E�5S�
�A8Ь����ԇ����:�����N��f���l��\�%����v�N����lb�yb���H��[�����1sy�t����D�#�9�Q6pc�M�� �z�iC��LTf�D�R���^_�S��G��~Ro��%)��0���)�B5L���@������*`�I@!�ǹ����-�|�1��bNF�={� �����j?����7�H�Q��B4aF]�o�>�f�xg�ʜ�}���� �9M�ٿM��ǰǁJ��̮�d>GQgQ�˴�:C��s��4�Q����}��ԏѠ��F�;���!�P6]�[�'�Gz+ʭ�ʂ9Y������}by-�'���4u���~4���u�����O�W�C�	��P��/6���a��諱�	��s�����i/�=�����)����|�W�Lo�2�eu�>`n���Y/@�ڭV�s�G`?p�uq�i�(]�%3E��δ̞�WS �qʩ��ٌ��=���ŠЦll;enOk��a����}��9Xm�9A7
�jt�Dp#��e721��b\Bk����{ZU���Ę"rW�Jk�vP�F�&����}�ĥ��-�P��91cA���:�R/:�q�4�;ĐBf��L�������ܛ�g1�����5b>�Z��IX���4Y?/. nD�l�Hg���\\�+���޶�����vf���(OO�B�YgM\���
J;v�b�@��~UqӫC����:P��a\��@<�HI�c`^~�� �$Z×C��\��2ʚ�Wm��7e��g�S+�s��?���FʒÁ���ƃ�?!����X�4�`��Ah��X��$�H r�<5�{���z�Q��m�nW���i9�(VN��*i��UYh����V�����H4L�LQ_h ۑ-�ڊ���R�d9�Tq-W>eze�.������T
�vas�}��P;�."�| Q�kg�'��i���k`�x�/��a��_{�����������~x;�XU�o�AW\Dn�F�ʶ�,T�=z�S<Ǥ����;���b�]�����T���v֣{��zzk�9)��[hY�Ղ-w�'\��`�K��ڇ�Hw���D�P'�H�C��H����!đ�J+6s�M�٨�t)��:f�i���d��H��D�J�ĉ�B�!<A�%�<_d��7�\T@����wrWw����d���iqަ�Wb�� �f e��c��c!I�v������p���̢�d�DDX|0{�9L��lE�� ,N|��d�|�~�?νܥ�뢰��������m*�[e�ow&����o�E�R8��H3��Yv6 ֓���D�:�(����TRn�\����>DN
z+?H��F�$��6����\�{��ɬ3�A,ɀ��s��Qi
�L���E��p"ٻ�ͬ�E�khQ� �6�i�U_��w&�E�{�����Y�dRS̥�������iT�i͋�К�sұ��?�t�/���B��O@P�k�`�E�N{���;��� ���3Y�8Ք&����rގ��mT��E�4Hd��ڿ�<�$�@mB�E�ƞ����R.Q`TG'�����k�bId�SM�Dz�n�9�I8H��j��T�+9B�:�5��5SJ����!�� Ų*o��q���6��*�X쁹���m#�����h2l\�������Ў�_L\e�!��}�g�j|Lc{�%�	��`�B%�I��-=�a}N���sj�248���FUU�R:q�U�+{�p��}��Q�C�JXWs�ٲ�Yۀ����b��Ғ���V<�rS!�a�M���#��
+<Z*X�z���z�U�mM8	6>��H�{'I�mp�υ�í����E�Ӄ@�G��"�~j ���ä��R9�4^���E�?~D�z��#�5����㢌E�VKuu�C�t�.0;k����]�(���E�caE�k���5����L�OIl���9������j�uB��wb���6���"���#���	��N��ծ>s�=�| ���?��<e���)�3x/���4a(r�fyֺG*,����:�Hy8�����}.9R�n�2Zy��B�H�r�_ l��e�U��d��NF-(�~چ�_9#�qF)u��i�i]v�޲t���2�ɀ\~q�W{l#_����v"Y�TeN���K���,<.��N��&aK�8�w9�eY�T����2�b��?��͈L�\�0t��w;E�0�)<=v5#b�?T4��-G� N�/�XX7�6m$;�s~#�S�z�[��RNB���ɴA:-����l�Z���c�K^1F��Ǟ����,"&З�M�z"C�*��`�CK�p�|$��'���k@S˒�t�Q���˚"�f�ngH�1�CAfz�L��N��x -��3��W�4.xm&1r��/"W[�DXc9���\IU�������]���XZ����u���������>�)��ā�Iݬ�����*F�ҋ��Qڃޖ͖J��R��o�y�E� �l�?�Ӄ��喇\�ȕq��Y1J�L�6!��uP�	3yU���,?��%����)\{��Dd�gI-�ݞ���/'k����.�
[���9��!,�3hf���oT�k���;45r�_�>�SA^�<mX�tݮ��m���"���U8���O��n\J\����4��BY���M��R )��{%��=�I	���t���Iǚ����n�8Ɲ�1��󍊹��^9��b���C)��ĬK��Z�0n>���O'Yd�1h������VI��2�w�$/���X�������r���q�`�<����	��a�p���t2��I5�z�[�Ė��jOV���sL+ãaeN���H�H�h̍��E{�p2�v ��]��/���ۯaVRiY�����/�Om���8JV�>z螢n���,H��|��>��q<��YU��b�rJ�ޥ_������y������:�e�(�I$$�~s��X��]�j5t�b�0�)��I�S��~�Bp�����	������&xUyO娛O� �sL����E��|d9:�߬��"?�)�-���{��@v"c��)��&2��?McX���e�L�h�,���ħ;꽜�~
�8>��-l� Y���n��M���v��^��~2
�Ɔ)����f�Ȋ��R#���J��uO�\�y�-	ۊ�ֵ>H��S�m�T����:��<��HK�Or@xX\A�7Q2JW>�5Hȑ���(\:���	S��X{�!����a͝1䝍�����g
��up��Q�"_�3��l�xp�h�RàS"1�3�lf�����f�%�!F_	�.]�Ü�
&Ev��"vO�l�1����=��Yː����x��uܴC�lZcUa�qAM$���/��"x��Y?��s�������[H����5Һ ��3pMv 9���0B��t�/�LNk͸vA6�����y�8ز�pߨ�ڒ�}��������S`{60:]c�>�{�~�f̒J�����d/г�z� Jz�~�����A������$,8Ø��f���� �ľ@����z\�°e�ofa�e��E\挄������@9b+[�4�P�jAQ"*��:�(u��\.�
�8@X��ʍo'�Wd>\��4�>A�l�!��a�q�e��;l��L��S����\��g�0�L<�`77v)KzQ�X�Sa��zZ����0;��8�9�����:���fA��"8�Z��"�5�(�u!Dp�c�iT]�ȹ�O�3,��m��׾��ǉ5�� ����hy�z)]�Or������@q\�=�k4U!A��}����E����R�v��#*�F*H���юd��8�	(�I�?�ܟ!E����V����3�~
jYFv�.T�ޭ�E��{Ǿw�NMI	���FW*�X';�m�i��[m'�X���{v���J���ȧQS��V��DWFf-��������K���~���O�2g��H����Aԥs2��/K�z����)���Zi9��i�wu��V���3�l�Db��@��]<���d�^��ɼE΄_W�(���=Ϡ롽� K�����F�V��?�9��#������fViL¸<S^c/�+-��g58���,��imv��>\3(йµ`����2Y���r��"a���p����c	lZ��/�on�(g��u�!(�4v��p&��������ݜ��w?�{�J-��i�`Y��B����)�Tڗow�]j]h��A8-N%+�.|�M��5�ӏ,t�����{�X/�+��,���t��P��t(�p�Ź.�����4+��e���BJ�Jv�-*��0ꈀ�ǯdײ�ċ�&��ܯ�:YN���e�S�|G}�����	�b)e�6�WW7��퇾��5��;���ќt?�j���l2��9� � $���b�o��:�7���/���(o.��]�o����5�Ȯ)�72އ��|�����@��C���
� ��Y*TZ�-�1�wޔXF���}]����/ ��y!�qV&�V�Y����M2�R���ȇ�b��:����+Ѵ��"6W���cc�p}�b��� �W�ɼV��{�b�+�� �lɦ�����j��db��M��3X{�>޽M��c7�u����_�K�s�I@�����T��I��X ϩ4�#��� ��v-�.��L,=*��t�;Ǐ&�շ���eLKH��.~<;.3w�<�.��r-Ho��Wۧ�"hE8��P5����6P9�Wj�!+?��d�ޑ�>4S��(���:�.$���
T$׭�Y(C1)�����`��HM���ڿ�	p�'�[�V���%v}~|(�ӭ���� �D�x�T�zBG�t
o�����e�Z)L݆�j_*���4)���i��ի�"��P�[�P��".��`gCyo�(��(��~#��,
�ySfH��Ϛ��+@�7H���
OtBX�1a��F��l�ȅ�r�x�f�M��2���2�0�x�ݹ��{��EFgl;/����k�%ȅe�r�6���۰́��#�S|��]QmqA���5�d����ly��{���ܚ�<LuZ�gw���r\����t*���uR�p��p�lㇳ�pH(Z��h�,]K��S=���2+u�[x�=������g���T��M:},�بBڝ�K%��1@K����r	�W�8F`U����S-J���Up}��x5�y�l�����;0Dz�1q�Qe9��n�'F�O���� �Z=!�[�cixT���=t��N#:�Q���:ue,��hK���l���D��lp���W�G;o��y4;)gzXV���۵O������j3�uq~��d2<����fؼY�e),�d@�:���P�J`@Ȗȟ崲�lJ!�=x�^Nv��km�$7�
��>���/����ݏ��-��d�i�< ��Q�u!���Z/)�u����ƃh���2Y���*c5H�1����c
F��
b���X_^@8<@vo/���Z��=!��e_�7�*;��񛝉 ��F㊾w�";O>�JqW��O�d��ts�9'���i�
��e7�+�T'KN��M/X�U��e�Mn��>]Z�ꩈ�$R��b�o�p>�2ݷp�l��bzP��/�������6���l��r��u��J����P�J����oaM����\��5�-������H�%g�ao�i�d-�C~���n9pY���s�_�=J^l�m����e<��-�l&dY� o�taЄ%�	Hn�P_�OG�+g�d�ϭ+h���.�|��%1�R��N�9ڕXc��y)�O���Y�oD�	���T��?D��nx��1C3,��?�����ҙ6���B��ٱ
q8A
~p��=�s ����� U` }ӵ(-�P"�K���2�~.��͡���>@$��i?)J=L���HkƢG�����u�%>�ɵ��¶[�O��"�4a}d3z����a�Y+=�)�&�:�sn�W��Éw�ڢ\��Ǳ�H�x���y f�hDql���h�?2@��bauw�L��8�KL�;?�$Ho�"��9��ԧx��<�ĊĶP F���F,y�c�|h�^O�w϶[�:G�]��׉�52�g�����h4Xޒ�YYץQ����0w	6�}.�Z�j�ſN����r���j��-b�pGH8��DA+�e&���nfBdA{����E�P����u� ��9�?*k&	=d�^'�8�B��rm��o��H�A�𿔫%W������O2 n�N�6|�Y�������]���)I�8S�/�����k�~>zE�+y��2�����[%d��?�[�r�FQ+�V�؇d���+x�U*H1T���V�)�X�,��?���kO���|��'ߎqk��X�y�#(���K��m��N|~�5��;��n���c����O���?���~�Qz�U�]��i��XL?�8�Q�x6�1�ɣU<��3�;��娜+��Fg�[���M϶�S`<� "u2Ei�-WQNཌྷ4�4,��)]��6�� c�
tT��(��{®`UL$��뼃`_��H`ߓ�ۋ��p��8�e��b��sFϴ�Q��3��#6+�O/�q�����$h����+RW��/Wr�DX�$��y��E�i���l�7'���ʂ���y��P���W4�Xu�{:�WERE}�&���tn�[>�$���,��Q���۲�=<B����c�%�5J�d.6��Sݕz�0�IN��7��#�a���7VKe(@����ι�<CȰgɠ��݁�Ӑ�3�8�aP�
<b� |�K�J�pm���ɛ���E��P��Fۥ.&W���_J%;Ͻ��ե$�W��4�iR.����٤|DZ��.͵��� �c���|B��i�$�[�jS!U-̰��w�Y�2��q�	�R(��j�!:����Y�O�Uk?�����I8�	^v��)���Q�z��~^P)d���Y$Mҷ���<�2�ٮt ��k�(�A���L�3@5����"��C�"I���x:x��#��~ޭ��Et[��!��Qյo�4���!�7�#�(�,HCч��׌�E�	�1��T����l��6I���m䐁j[$�� ~2X�ip˵\�J=��
��2�T9&b�ֲ�2`�v4�0�t��Ҧd�D�3����Ŷ�=�y�&5�׏]��͂+ Sʱ���e��0|�b�H �A�H��1��%d����U6 �IΒ��0,���iRYq'ܝN�! �gz���,��H,����&V�ozJ�M6�|Ets��>/�wMM`��1�?�.���L�P��4SQ����7�����O|P���^e�.he�@{���Ϙ'�=�,�2��D҂��a��F��2!����!���BR�O��� g���[D��1g8�5�s�m��PH��
��;b��<�.n�8�"�9Ü+�#Z�n��j:���x9�y_Z��Ui&��Zc���T(3�)�Q���u��y����?XGU�7��7��WR��F��^(�Oف���v���ۗ�x�7�� <�xWn�rh��UK��n���+���_���6�o%��!:�cb� �Q�5����zX�V���qoɶ�=�s)I{��i�L�ʋWS0�-F��R��~��r`W�_	NC��-��@0��",�%�w$���h(P�=
u�H� 'Qΐ���H�����Br��s#�g��^B�������s�Z��ҝ�Jn��E�K.�z�bsBo�B>�^�E}�YPAF�s���t���d%*��"�����V>�q� 0��o�:�β�Ŀ#�U����M��nE� ����~�+q��$����(����/W[
��t]է�x���$�Хz����e�:�_�)w�Q?���|ϻɵQ��7������z�_FJW�$D���"N��K�S��#�0��������?�C�=�pO�=��_��G��Z�+�`ظ"-��ZS��'�%����R�l������;�2B�g����:����rz��5�bwf�q߄zX�ΟsF7
�]2�~��J,G@�� �I��T��R������$�q����!�\�	rjfA�y�6_���R���?\�،d�C�ɳ�F}K(���L�����j�-��|m8�=v�c�Jx�A�y#��B_� N���?���n����]�Ջx��M����k�X?�t(C�<��h��qyG��ћ�0���{R";r��D�B�J��|9��o��,��4�����(��PCsE�U���샴�%uo�VW1]vv����m��=�@�k�61���p��*�mq ���An\n�>�>��w�P���Р�I'�Hɍ��uz\���Σ�_��9�.J�it�'>�-{Gv�l1fs���UzS�W�N�>�4oС���1��P�Y�[�a��|<8c�`�V����:<g�ZG��d�U RK�m���J��}}Oy�a`�L���'0�T��X�	q )%��r-܏P���'�E�g;���)˪Y\�ڿ�g�--m�2o�5�B
�r�*9;��7�ٻs�?=�W/h��J!�C>\7���1� nSm>�A�	6�/v���^(�gHI�e�^��6�X�ݗ�"�L������FQk�N�
{��w�[[��L������+B�h�7蓆Bո��>�,Lχ���!P���'���66o�[�(�Ni��w	����F�Bԁ$Lj��9�jn��Y�)���i��v��23y�Y�c�o�Lo���L��З����a̟�1/�*���D��B÷.LGgv����]�n�&Nl�$�}8�!�Kpy���q�C��)����_h?!=�V*Oޚ�����F�^��]h���+�J����#1e�>��Pl��O6����p E��c��\���XF���(���f؍Ԓ�z<�"� ��~�C�j=�J&�^M��#d&���ʜȽ��8m]k"Ȁ]��R�Ed=���D���V�L:I�6������|":0B�T�����0�7�g�Ư��}<6���c��%�� ���,�:=BoעX�$�K��>�"͜lWG뇞��j>cا�yқ�LAM~p��V	�?l�m��b�
���d����ϵ�/5��
�6q���-��3WC0�W��S�T�*R���k�{R�Q�,Gt�wh�&��tc�2c�̴�o̓zN�g�nܷ��[�"5�Tw�=O�+�瑼MB��z�����<Ϲ��	G��2��pl���2��M	�a\_�3�gL�vK��hR��#P��ǟ]Cl���5�gܒ�U\$�H}rT-�kᑜ���CJ���*>�w���/wgp
; a�:���.����'r�c��[����u�a%q.N��1�?� ش�]�*溶�}�kR��{��֜g���\ÛϨ�q���Y�S�JG�I �*���R�#����&�i�鑒�%�ꃐݡ#_�<�1x�m#�H�ZNo�w#?dw���U��x���V�jX�&�.�͟#�6�XΘ�~OZ�d� �QAG�w�P-���}ܝ�w�����U2��yax621����'��O���!�5�g�T���N^/�����ڪ������
��ډ�T�4T�uj�m�����䄖��
p�c��l�m���E��k����,�l�kؽ�-~"pB�:.�ȳX1���|?O����o�-��П���	�������  ���{C��@��V��7| �y%k��5(�y�>��"٭[��ۮ��^�'��@Zꦞ[�-�N"�K Ψc��Q3�c��Ţ<*�t�h@�'�v`�`Ɲ֟�`BT��ec�W�r��:"��9Q3�s���.��gg4*e�w���4�����1j���i���8���-�DW5ҦL�~��3ʧ%E�$�AFJ�9�MlH�|��Y�r���+Z��w�s�|\�V��'���՞3�g�؎��з�E;;.y`T`(�#^7�5n�n0��Lpy�����j�(O؎|�n��Ds4���jD��2 ��?}�MP�;Z���i~o�R�rT;k���������y��;��@e�)�A��.R2`�ҫ( %����p��gp�a�)�Y���W���2�����יᒈ�l=��Lߡk���(w��N�1���[�;o>\�����Kc���5w�3s��X+����ş�@SMd�k=9(#Г��kBۤ/@��O ����,�d'�(��x�5�#�FxY�~7E���SL��Tߎ�[��>��;$�Y��kp60�s����0=��Ru�}F����Q����Ω�� 4����c)w��q���K��?���*5I�"ЬA
:X�2T��S6r��Z3z\�)˄���K��s�WN�[�<�ӢC��� ,�K��;�b��ںRw�m��A�լ��pww)���Kp�zXv'���*13��ʟf�z7�C'�����ǰ�+lOt��^=���"�=��ɧV�u�ZK|^+�5^#\Bu�y_-&i�j"�@ȟ�O���?�uq������/����d�j��Tx+k?�<�@Z����pfzX;�Aj�2�k<I�"�ڃ͊6��7=:�:�Њ�l:e����.D���;�C�]iQ�¿ZS��$����pL]Rk�\/O6
�R�wӶU�re�ӽ���`$p�p�=��M� ���ࠞ�Xԕ&+�F(`y��~��f���y�Ҙ�p�j�0�S�����0��=�0��Ӗ�@�2��eCg��t��O������e0%�OT��t����}I�!V�"#@�Zн�-�>g�ə��]�2�֩������֘{�K��)�q,l�N���F�%U$�"�:�j+�t��o��	/u6A��r]��ܐF�/]��й��@�!X�U�g8���� >��&#������B��M1P��s!HZ_�T�.��k�](0�"`�����=��"�ǖ%�7�42���sܕ�qj��<���q(��k�5�'DZk��3,���3��ūo����*��8BGN�B7�Beӹ
��6�2���*g����c��*_�����ϧ��19}�z�����O�Pe�A��a��>��
q-�r{�x�,
r����-�r6� ����-��]�c�{�k���V�>�#;Q�j���n��;c�������Z���������DX��1橂+uY&���n4��Ըܶ����z�pDT*��89�,3�,��� .F~�d5<�������/��q�(O��Fm@��K��^yh F���#��3-�|;ЪJNߣ����|%F�$a^Ҿ����zIw�t�	���{�g[ߐ|��>0D�(��dʑ!/4���c�Jޓ��Ç�m�c�M�}O>J��]St�vs���l�aa!��}P�e;u|��cSː;*ncP�K�Y��v���oJ*H�n�yנ������Qܠ�)������-�2��ɖeH�,��W��"���?<�#���
���4�B��9��B)W��3�k8 J���,r�a-���ܘ�n��)ɻqz�N5r����W3�U������b�r�I�A[����חU�QJR`����mwQ H�$�EBg[���"?�*�
?#(�(m ���k�X�� ���!va��y��C�g���t\$2�a|G�j�P���E��G�zBf��>̊�y�+��!h�.��G32���3���;��7�잷"s��X���i�K
͜�:�F����s�wY`�Y�6�ݺ���|��z �L��,�0	0M��v)���2P��ăg�I
憬��2'�p���mn�Y>�4Rao�sp�����Ԉ�NOi���)]�^#��G��m����D	.͉M	��]8��#2��s po��u<Jw�f)����z*�a�)������a�}���a��2i:]�ɗ B
��[8�G�-aƓ��GV�R4��]@'/
��O��	�M�XJ?�v4�i���\�����gX��U�����ٝ� ���Bq_xO����KA�����2?*�2�-%K��bf���0��������a\��oǪGDW��:���i���k�B.�
�I\b=xl ��X����d�<���wp���� vi`ԃ7����7Iő��C5��=�`��|Y٩��W�|�E"P���+DeR1�<�w��p�r^[cNc����hN\���?9���̰�?���٦�oj�<AwL�Ǯ�S���x�$w�!���x'VB�e��،=%���0���*��);-3����/�99��T�d(�h����6O�#�V��R�W��ohX^����:�"Ɵ	VT�_� +���	�����j�����TV��;D�r��1�e$k����'��ôkU�O�M�Oĕ}$Q�r��<v��,��E�o�o��� �¸M�V���;��P��4���z�6�8L����a>��mU�n%��ej�2g��p(�ƕ��V��򦘸�_��ψ�t��q�+J�>��\5�n*5y��퉇D�1m�'�/���vR��fч�K�s$<��6�mJ�s�ƣ��\ً@��7=�Gp ���+�����{��-�.N�Q�����)���,f?�ҥlP�E���>�{+Q�v�.�`u���]��Ƃ�_��	�oխ@ ��C�"BOӑ��K�)�}�{�x^.�������y�M�rW�֒ZX"��j��^�6�."�姉Zx;���fy�i�5z8){j�i^'NG®�Bl��h:/|��������1z�9n�B�z�8�Vr�h:]D7r�
A(C
�0c!����J��`'�|�����cf�眓�*y ������y;�;'	�߾�)"�q�,u�u���7��e�!�n׆E ��>&椠�^��� �;��3�7�u(�c{6�U�j?�L;�叐���I��yг�>��i��vdث�*|l��?�x%ID�)��KZ�͑�k;�.�iZ,������W����L6�s�!u�bgk��H���K
��0OUe��cх"�j�"�n�
k�{�r4�2b�z�)q9N�#g�-b��6;�x(�05%,8�y&�0:6L�N�?)�@�rc��?��!�!�]4�J	G����w���iX�M�zI<�}iS�d/����E⏐��v�T磝� ��GQ��A�	�w�^��q6��c)[Cz�1�H�O���>h�m��V��-���#���8����u6�n������@a����O��s��[x�C�UY�����S�~4X��3��ݎ;mJ;��5���?��*q8��[�P4r�<ܧ�����B��Ƥ�Hcu�Y� �J}v�3��])�y6����{Ӎ 5�J�ID���M��+�k�`Ӹ��G��`�+f��^\�������a���n)��ô��.L�� �?��P���P�_���I�!��R���W�A�)���(��&���9��W �iq�w�	t�n������'�hy3��D4���N���w����Ui������h��Lp`�����#�RC>?�����=;���1xN�m�J�]������o��w���&g1�������n��a@Gn!	2�S|(��Q�ʫ��7���g�d����o�ز��J�Mv��@
�q�pDbǧn5��q�\�@�>ॠ���'�I1 �	���Xlu��#�'��V��iB�uXd��u38qGq��,���Ӧ-ˁ"�r*�����]j�G�.m(N��D����l���)dj�?�[j(7q�:Z��J�jP��GRϫr�[�2	l)[G�!�'1��2L�D�^a2u�7��:2�B�����&X����;_���'�'��Gd��W����`6��%���,2>��?�����4~so	�А��^� ȇ�0��3���i!��ٰ�x]使;����U}��3&1'����1ȭ����V�Y����[a�&�ym-U@/aZQ�e�d�[ٔf$pY�Ѫy�l��@w��u�Ӛ��>������] ha,U#��Z��������4�Y��9� �5Ρ���?7�$u����:Lk��v�A�������\_[��S&�$аH�a���rNB���$�	,�T���mX[e7��
N�!U�0�tz3Is�w2	-t؈�YXO�(�`o�6�d���F�t�l7K'#���j��m����%���������2�EϦ�e�~��`v��rJb��Gl�\�um7�_��K� NJ�V��.P���{O�T�Ny����}�a�]ҵ�V2=�$Cچ��nPoɵjJ�T_.�U�*��z�*~ꯒ>=r�8�0���_K���q�����^C���|���nv����?cĽ!��Vڍ@�EB��5���(�UsjP4���)���(Խ�\
0� ��oL3r얮 ���d܇i�Sū�"��v{�=�t*�%�Y6n1Z.��𛳇�y��.p�|bE�����쉽��_2��Q4�=���j�V� e��Ir��yb��	�{���^��ك$�ɯ��Z.��#�����QP����a���e@Z���U��^�tR��Ƌ#�q��l�l�}~d�h�}��o��iB�������fu�C�Wۓ���󤀾�X�ā������/�'5{���,U���vcC���@�m*�O���E�7�WXj3���齩����Oh����4��޾z��Q`f86\��a�L����q��eϣRqT6�Lu(E w&�"7�Zm���72��0��G�7p9�A���^4�xn1?f6�h��ޓ`q���f�\��
&����|k5�x��R5 
�2�ۥ;����ά�� ��T����p�\�^�� ��_��͂3����QA�5�h4te�+�I�x��|�c_��l)ed����  ��Ho��?����x9g��v�Wv����+_�E��f}�}��{i��i�����$�T\��ݛ����?��P_V��ۛ�����*&��!y�ً�xr�}1߅5��q�ѹ:���IY��&�ާ��zl�����ϝ�v��ۺ�č�I���JdG�$��H��,�y��·�/�y���r@�����1ܿ��O������Ħ$�E`�)Ka��W7~.=<﷌�}?�j�X�z�!������/ ѽ9��p��[�QSx�jy���%TU(�~�m�����Q�|L���Ǜ��d��X'j+9{��i���eO����������@	F����:uQtpT�1���ŏ�p8]�e����=}�m��*���	a�Vd���`��&쪌�<��y�����֠�J�c�<XDbK!f�S!VLl����Q��>�;K��~!GO��3'��]|������
?��͕��ԥ��_��VR��� +�|܊���^V�y|��N$�@"���Ԥ!�&|�s�$��p�a���v�;k�wU$��ͫ:��0b!��$D�\ c�L�I ��ͭ��X���S �L᚟C�5e��o�J}�o��-���{���~%Af���Z�Ǝ���+!j>����§j,�Km$�Ř@D����:ߑ�{�x����Mʱ-�=��9�O�Q�
`1=��>�ԁ2	��2�cf�A�AN����P1��	(�~*ו:5�1��8o�H�:��"�bL��ٰy�0:�^,ޘ�̒J�&������9Ó�}!^��j`�9���j��X�*���(�S�����Y������&��/��A���7J�:����rRr@<��)���kr&Ȅ��=�N����N���~��YG)~~~�ii�x*9avc�MTV]̠�y�d	�a�kgF|�18�q��|��2R�� �QU��Kn+�	��^d;_��Jav�2��2G�
5FGC�B�!D�& ~���磩�RV���Zf�j�L�/l=������ x���r���X3�c=��IO^�s�O����,�}!ߴ�&��,�6�*���
 o�h���uC�>�w��_�{5�
�~ՄgU8!�aQ ro͎��n�\������+���b�(�[L���2�WV��!��rfˀ��Q6�`N��4�)�xDOuL���#-�?H������a����JG���C�X���p�Xg�H�!�~��fR���H��/�b���>s���?� )P�~N(؏�+��$�OX9��������Q�eS�
�5ۈ��e�3���^��,�uH��Z�@J�K�ϵ�V1�1��Ŀ*��8{0�';�l6�I���S�AB�����R��+W�c�M�h��rI;b�4ɣ��E�uS�4�೐*<C�oֵْg-yֱ���~n^�\�-Z�������z���7�(s�6"�E��%5SQ���Ă]��X)���S;�@��M�ti�#��NA�55ܝo�fM&�|' �^<�)G=�u�^�F���!2��P��:�«j�@����W�Z�cs�iYb %���H]u%43�}���b�ߤ�.dMG���4�齮N$v�a������@�u^r�g�����E��t���L,���xu�CK����u��C���=����Q=�����5a1w)��:�z|�+�QwN��v�1<qvd�n����Ql���>z"��?%a��Es��Z|��b�hD�|�:�����|[���v|S���k�v3	w��>�,=�p~w �{�h9!���)�A�%&��
���� c���% �a��6x
9ꍤt�95nA|��2+o�E��=��>-pk&.69?Q�>u�[�R"]�g����Z,�5 Pf�M5�c0� T�b��,`�Wy�>!59�2�8�BD�p�iB*	�\ɨ���,�M��~P)��#&�:N����W^��r�S��L�Y��NF�Γ�@�8�^���؁θ������,n�F+����Ì���p�<;]Gs����Q-޼3�⼐�C5���)��Ǭ�չh! l��'��>M;�.�l�=R���Hsx�%���PRY�ZH������:�˦O�|PP;�\�i�9�ZU3U<��Z�k����Xl3n�,ąf�p\�N(1"k��*.����-�s:8�obX��s�n�Y5
�#���,����O�"��G�o|���9�#i��1��Z-��2�XҼ(7D�,�N�*�c(����� ��[� �|���e�Ky�d�SIs��%��091�#����8�K�������L#���4���ڒc&׊��
6>��co/͆߷���@ŗ�|���R��鱧*�(��^ ����*����zG%������Tu]�3哫s�i�Y��/.n���V>;�S�N��Ly�lTs@5�fa;t�����N�!����4H�㼤�,1��nL�����KЎ�ڲ��_N*�1P� ��emW�.cT�+'=q&c��T��65�~��}h�,_��}s���/��U����)$�=պb�q��2jW=��"�F�Hee�s��Q:5GaȠV g�)Oq��Ң�$��az�,^�%~�ʤ۹�N�3m�.��vP�3�K�ׇ�}��<t,���1��F�Ĕj
�"p7H��-L���c>����ӽZC�g�B���Ĕ&��
�K�`5mh���M�-��-A`a��篮�5��I��wV:�	�:�0�e�ڒ��k��8��<)� bt�x�xzM���P��an:)�agrrii���$��h�䂓�!�,�b���
}��Icb���ߜq=MN�'�.�9Ѯ��[����,��R A�Ӭ�����y�?~JO`R���7� �]�z��_��-ţ;�(��C����~5YJ�&*�jp�����M!�00v-ř7���ˁܳ[��:�F��G��A�aD�n%�r�h�E@���}��D�g�H��r�?����n�<w�W�{t�3�}�T/cnEj�7:�HWٳa��[�-F=t��X)���E&�6U���{��cm�d��G	�)U�aD���F�x{�:ұ��r���C�����^��!/5�n4Ԡ��D�6�5������TX �{J�]�M��!���`�})�Ln�@�k&�|�-���+6/��$o��T&�[�����@ɒ2Tf  ��>Ƕ+�k�|5X]ض�!݃��q����F�͍��P�ݹ�"P�CyE�"˰,����d$�H��{��A�GqPκ�g�w16ಃ��(����!"�h�	?�O�eG�%�{n`��F�2�����4]G����NB9�ξ��=�D�B��^�%zWAV
�k4���B3V�0ќ��D�\�6�Z���^�%{<G	�A�|f	O�M���������5� z��t+��ݘ��t��Y ���8�$��2.E�i����<�gRȫ63�C����\�I�2�Cc��i!l%L�#���Ѕ�	�"Qx�2&U`ӣ�Y�^ƣ*kܪ��L_����XC:s'���%�/�~$��)q ���ʤwx\v��Ӻ�t�݈�txr�����y�Pz�+@�qD��ێļ�����VA,.��*1�ZQ���-����B�
]�ƣ:0�'n�i����o�@��_�nˡi��څK�3�����d/�� �������ێ�=�.��7sB"����+0�u��or���^[����\!�ԩ�2�s���
��+��� ��&��5�q`1N�$��z�w�\eaR���#ܩ�qL�6|�����s�e%:�����AG0�%���8���Vh��W���(�d��(�g:Ŕ�d���I�@o��\N�}`<�to�T%K	
�\.ɒ�M�bop��Dl���H(w��#0Hݔv2����U/J[(�\�r:�۟Q������h�K �)ym^ON��9k��t'��u�~�޺��F�vz����������C�ɪU�>F���$G#	�M��Ɓ4���c��N+���t����1l	��snDkAV�|6��E��IK�������)�����U���Qz�c�bo�d#��"�d�LT�}̋S�&荋1Z�uuAV�.V��NFd)\�5��C荻KH�,�?��z��?=��Y�]ҹbى���(7mW�LL�]��@�N|��\J�.f�j��[�4V�X�9�Q��A��㝵7Ƴ��mcB cg ���C�H�>��*V��}��@s8��a�QYm�������ʫ���p&���Tk]��y	$�I��tP�Ψ�A��b���J�*E	RP��5i��X���mW3�嗯��aZp���X����m����2v�!��;��7hLn����.=u�gg��%x��E-i�;�$uRy\)�_ :�ou�/�g����]��R�'%��U�t�M��2}+̗81vn��,��_�� �;h�#��q�r�n��\�"��ܞ�<^�N��N���ܨ����ro[�
0���*�&�^���Z���פmT3���"qvƓǘ�˘�[���d��< �:����}�+�A��\Uc(�4"C�Zlw��3J���E<��;P�No*wv$ݜ���>�˥�&�x�P\��X7-��m ��ծ�'iz�'�v�����b)����V_�b�'y�-���(i���1��+��OL%Y����^���^�׃L�d_M�b��:���^���Hޠ��Us�m'm}��hO>��O�`�k���*t�H��bO���1Y��!u�?~�GmFn_������f�(|�Dk!y�R��%.��L5zhe��lDYEyt���r�@,����=8��:c���j]��&p��?YWK��X�
��'l,�r��Y���Q��ˬ��*��9З��h�ٓ��h1�ni7I��k���4�Do�8x�vy���� ��s��%�!�����T�iT������c��;~DZp/h�"W�Q�k�<�(W��PET�Ĉ�H�E�4k��g,�:�8+��?���=Y�~V��pG�Q�b;��	M!,�&&Y���F80����&�Y�Mm�H�,��t#����;AY7�5����'�%`p0�p\TL�/���9��w��܌����@�#䤓{�Q�>	���ojwg�ɩ� س2@��w�?˷�XS�m5��{H�@���Թ���^��Y�)��oZYH�L�|:;��R�"�k�cR6��+��ikE��	;�h��e�o>Ok�[$�\�b���T�8ZȐ0ﵨ�p�+ę4M�xL�%@�;/�=C �qރ�
�3��N�c���|�;�s�L�Z�I�_Ȩ����E8mOH��-L/�?߹��c@�<_g����\��&�5p�e���(w'��*��Sݞ�h�rH�S����*"�0wBr��Fq���7�Ÿ�k.PH��>;�^�^�V�k��F�2c__D�3|�=�*Ý+9����$�V�3�����1��aG���2���5Ao�GY��=@󦧆'.�p��D�\k���
ץ]����}���ȯ}�&a��x�I����'_@��ݟ-g�ۢEn�x��%�ײ<�nF\DG�<]P�o B���: N��IHl8���n1M�[3���ִ�=��>���R��R�;�	C�d��ͣ��`�(/F.ph��U�?#�=PBa)��h:�j1iI����Z{���N�-I��l�R]�4������bU�nѺY!v/Ե�r�L�y�:a�؏WV~��UZd���jR՚���6@�K�y:�����0��t^J�� ң��S��e�ez��k.2hT�@�|Ot?�ʈ�.��*ۙ�����6Q�f n�����LjL��02���n���:�0�FE�ݍ���1Awy���21�mu��7M>s�#��*4�)�z�4~�����P6P.�`	�r`L�ĵ$(���	iF~�$V�D!A�
wYɑh��GE�7��^�-iZ��K>������O��`�)M?Y������)ָM֖�3�o���=;D���}����ؑ�sh^��
=��щ6�m�7r��6- b,�<�a��d�~�3���lR�@�_1�#�1J�7�A*n�R�d��͹��z�I&&�ET9�X�Q�x�r�zy�~��o��(�ڗ?���l�?�f��I�9/�E8���͂į���]n=넙�y[��f�F��)ܒ9��y�����g��F���mO��iΑ"�0b��� M���Ӓ���;�=�P��d�?�kI}B\�[L29�%֖s�q��iR6o�+%~��X��׼������í"�w�n�إ����K�9(*O4B�fmˆ�A�!����
�)@viN1�m�.D��fl��9i�P���Y����9@
���\a �V�ݞ]��-uoZ5��3���$���?�V֦8�/�Ma򴮹����l����
k�Z��g/h�ج��S�Z�NC1MfR�":�7�rE���%x��� �����L���<����?� �c	G���~�AP�$
~����Trz�k@�9ЕT!r����FB�X^����Z��%�3��)���翠���ޟ]���;�/���Tx��)e:sV�9`��gF�V���4�ݭ)Ak�M��Fg��+�I"�%���[�|���4,���j����<9n�D���68%y5?��
VG��6��o,����?�"�]H�,�B��4体�@P�^9"���?�*�w6}I��ĵVBN&x�e|�1�CFYo����LQ���]�(��tCˮ�ۥ�����@�h-���ұb�jmhE��_��T�Ҍ��i�*f.�τ��V+}w��;�~D޾nWC9�àyheQ�j��m3osQ�!���Z���Hs���P̆u�L��Y�U:����YQ6��V\��iB>Z�L�h�5���P���Q7M<�I\�hk����K���]�>l��0�2��T�hk1>�I�]����	�*7�I�����`5�_)N���=SYU[�C��P��б�Q17�%]�n�l�~�o?�~���`�5_�`� |���6^/F~K;�0t0��s!R�o��f)
���t^,@��:��]��/4�dw��C(` I$oQ��΄S˕�H����6M��DΞ�S��Nk��lvmx�3�k*�/y�4�v�(%m}�i�����d��.����ƿ�qE�����	_s���U�*�������ʚҩDAP�W�/ǆ��`��籵���$6��.SY\Ӿمm��{�܄��1:�mQx�^��FO��B�ڃ6��tZ����7_ua��w�Z݊��m���U(YOC1J�w���V,�c�4���+�ѥ��U���R��v`Z�DcTl�@D�a��\S�:|�i���$;h_��| ���>�?�._��U����jIm���u�u���Nx����`[Rf��\�B�뜊<�iX��Uۉ�������s�����$s��G?��E��A�"(���J"Y�O{bY%@$=�=���unM�g%3>}2b��b~ D���r�-��@ 6G]<~��Hw�+E��f	��
-Y��DS'�4c����̈��+��_�
�����E��mX�[�tE�����<�$JI�L����\���Z4r��D�֟�Lw��p�poɹɠM��TJ� h��m�e5��8�<�7q�EJV-������(�Ws�[߁$��Fų�/:f��G/���j��x��ySq�V�C}(򂢢h�������F�9'��	��I����o~�e1�FQl�
��8l.�B��Վ�2 %�eh�S�qν������w�
��P0���va��%�X3�+�L��D4xz�h]!׷��;z��6��e��.(g��]Y���E�?�+-D�Od�%���S�i��D{����dh7�6�J<$\�k�OB	��CP#c�1!�J_�� �/J���n�|��
�E�igV-��M՚��zʅ���UgEӣ�<�s������ޭ֫�*氮lw��R~�(�Ao���,�%nîp��F�G���6jا����&8<�c���{� '؃�E2 v���V�.���Y�ۺR���z�*P�+2�=�� �E�T�c��>��uZ�y ��="Fg;�͝��Hjg��(W�Ɋ�͎���|���~�rLO|��IF��o�*G�dە��x�9�{k44��!/��!Ps�������=O�I�gc7�]2C(y��x�Gq'�iνBM�x�#o���ց���/q- ���@��,�7y?F�5�S*�\�� ��R���d��S���m�������8�[QCg��B�х���j�X_��UkFoұ��-í����o�a8�T%��u�mF�9ƚsZ;�`b�L	�[#/��p��-��<$Q4G��va�s�_�����&��$b�;�	��x�v�)2AVL+�㐅׫^�s�[X̾�.���V��?q���2�'|��} 8ĳ�����_���1$�.u�x�Lx:?�_�+Е�j�Zs��z�]��=r�R�tb4E-D�<�	��v�=dH�f��X'�5����H����w���kB�b@�+���jf �$�A�1w}�M7�_���<s.�-r����ߞ�Í���b��|'��䋷QAdi��h�%��e��Y>����rVfm&r�F/�o|eN�x�َ��r��1��3|���}Cߩ�s��bL��+��7��y��j�l�%���cU��bY�<r�?�	.�y��8G\��0�	�D��7��.�W�˨��%E ��ܛD��5Kԛj;ҝ�p����&Y�N����s�]�۹�лٿ;�וO���	�w��R�[L��z�[�� �ԗ5��"V�%�_�HA��4����ѓ*v!��,E���4��[nV-��Z������z�Cm��MzT�@���
-�l�C*�4��DR��9#Y����q�5�2g"&��n��?ɏ�1Ɩ��#Cܐ��b���l:z?)X������ު�F&p����Æ��v�Êsu�ڍ@	���p{����>�yy�VϺ)���44R�o���q� <��Ѻ7����ۣ�.�Qҳn%��|���`��V	{�U�9�6��P���s%�r���{�1�[h�_ |&]|;�\�}��t]�_E';�	:u����sF����/6	@g�u1dY�25��mPg�u�5�8�oH���
(Ԫ �;E�:��t���I�W�;����Ӽ>�cک�Y��,��$�/TP��"`R�1s���KI�y|��]��g�ik�/��a��ñ�{W���V���p�����B�&/��p�|��Y��v�J�;Un�E��aӞ�e��ٽ�Fψ*YQ\%|�7���]����Wu�e���D,t�@�%p�c|���+k���C|H�UG����=}���������A�5_\���@ ,f���Tb�h�;�� ��J)���d���%zI��!/���=R&�����T�b�-iA�8�%�ǿY\q����ie1߃�OJ)��S��Q�\���X޶;�GK,+�ߧ�����%q��Ӯ�i^1���.�F�NuWL��{�xn$V��c-0�?���1Q G!�((�"*}��d�Bʺ��h��$6���@R�k��x=�z�jץUzX��t�;��uV�<���x�Rk���,�*\5��s�.+�cj�{�3���nlнMȊ���yK X��KFO�z��	�4���y.�6� \h��Hr��>�J��"Q��\��[2��(����~��?'Ξ�����P�U*�P�a�`qGZypuH_�(O��@���q
�����pM�w��P����n/<̲A��B���MZxfTK++s��Ov,E}ӊs��ӓ��=A�$O��{���?o�E�`N��,�j޻Q"������a�� ϜL�>�+泾p��)��|wX��i��ibrvlV=�8�Q��T�~,ᰐH5�@&T��7Db���=�m�S�m����=�/�s� ��<֟ս4L�у24u�f.�OҞ�1&�:-1E:��!8Mm��q��*H\��Q ��F�:ۚ���X��JN�T}�ߕm7p�12�j櫇��rF�{�\��: �??�3ͪ����pM����|�����#C���D{��0���z=��Z�8"��^���ʻ�����Y㌠��İ(F�'G\�)�>9H�L⭮����n�^�)
�"q:����{F�8�n�T�D�#��ڿ��,AF��-���V��l��	����O���pD�V�>U��Ct��o���G+���h!�#X{�Yz��M'���l��A�?��z��h:̯lN^�dhp*�9�]�Y�� V��p�~fu,ޑ�3�xL�+�zƟ��f�4�5����h���VaN!����HN7<�,&1Z���u�a���9�Ձ��H��/]:"�;�?�ʲ�*@�U����Kc��x��ШBJ�T
��_��2�]|��Fǀ\�')PU�,kL��ٿ��,H�s�H�)�ݠ*=��	N�2�h��H �����!U��1��� �˞e���̋]��*��Pܼ�Fo������2�i=g��$��8����/^�$�t�=���7	�6@��r���֥79�T�Jῠ�׭��[�*7iZ|��9W���ي�W#Wz�����B��Yc\�Xi��1_���#Ss���̩a�N�W�_�6;Z���2ɿ����I>�w�(�h%p��	'"��5n�R%�}٢L�H�V"D6V1�x������
�{��koy��byD۩:�m�\f��7j��`OU�,Ⳉc��yN.e��e�5o�EC� �)G�,O�Sg�$��J�d�&4z��\��D�n,�L��5��������C+|la�8�#i��?b�K�%�c������E�V�Ùe�j�?�><�z��k�@�}����lt5�G��¦�Y�cF��&~��xc
aSWA&` ��"C)������<����mygO��@�L������#��$qI���m;/�71�K�R4����E����U�~*��F��m�u�l����h7�P�8xj���=������q�!yb��)����hm�p�<q���t`���j�e�>阮��U�nt�syw��k��>Î� �`K�y��3����j�:�;����[RE��2vM�*}ܱ6ñ`a�K�?Ј��
MҦ"n��E��ŏ}	σm��(��o7Uł��fd��?�}�Or��o���.>aS�����I�>zȾ�A]12��B<0҅�R�k���S�
l]�A�X���/P{���q�b�銗��}��!�t��L_�
�%���G�F���U6�e�0�N�y��z�ˑX�c��'��𕛥9��Ģ�H ��y��W���Mւ�r�ӢV�����9�4L��,g��S��J�i�0�c!�-�%�̡���u��M�>�qL������1�F����A�C���� >�UA�-;h��8\	�q�����͗Cሷ�����f�\�]��ġE�[���ފEq�!N�n������ >�˲����N� �!_WM��w3���W0�b�ݕ�-R�&��d�3֔����.!�r���?[�0qyY��3��;�KS>$�-��z6���g��R��%�-m���Ef���P��K4�I��b���J�[��w��7���q=ě|LMe
�ݙ��#A���{}pظ���W{�EdNps��#e�c�q���e�=��)y�c�eO�q�6H�d*�R����H�]���K�vnn���GwL6D��m�b��F��g�JĊ{n��V�
KO^j�ZYZ2ܗd�����\L97أ�=J��v�
�Y~�AbX�u:&��g�dcngp�Vl)Ŀ �s�Ӽ�_�2
�a,���Y��OSs�v�+���}��Kgyb����Z��  �3s��ߍs�O�d�f���-A9��7q��O!D��]̜�轰��5)S�
����%KFF����@;�!U�����(�ݛ���G����^���լ�p��j��ZIO�`$t�$Њו����1�[�4�����,+ba������ts����x�/a�������~|�oc�D�{|�1a�4��}k�W�cȧ'f�~Hz�UgC�|�W�y�9N ���0��Ϥ��لVR"v�'� ,9Z��`^~�IJ�Rp��D�8p��h\���(׏�{�����S[��?Wēɔ��B�)Ҫ��AP���.Z'�'�Դ�y��Ϥ܁�U>,�;hZ��+�T�k�O����(�O��AB���oE�ľ}�r� ���C������87���+@#�~#���FŞ/�.FFI������^ko�� ]���R�B5�5 �~?]�g �:�:���90���S��p*��}��9y�+Քa��_�~UY^fP�����Ղ���cI����l����Sl�����)��֪�������Gl�o�fauK�Ŭvς��j�������Ǔ8��gPh!�����8������T�
��;�NM�%ԛ��_m������ �YwG�SB�C���E^��/ GϜ�(J>� @w�P0IF�Mǡ끫�(�K���o䱲�{��a�H�v�\����9���ë��P��i'�7���"����n��F?s����5`XG�~� �IT�Ȭ9[d���VS���/����ޛ�i�)�>>���K���	�a�ʟ�s�ug��v�X��e,�ͅ��� �\�נ���+�R��'0����4�F�_����K�埡`9t�չ�׬0 /AڃtO������QGe��.�`RP?�`Q)��Q'��	Gy#%V2ݔt��培�!�䄂YW� g��T��	+��#�!�ԍaǕ#fN
�LO�ek������?����~ߙ��
�FV3:�ur�Q�V�kQ@a���3
���<�0/��=mX�$�	��%D�n0Wi��5c�^�k�5,G�G��L�ܴ��<��(h{+�/c�z����R�dϧ�n0ϝ�Xo߆�f�q����sf��)ˌP�� �F�	�(a�&Z��=+ȼ�������� m����V����\;��
�Y	J�,:t�4�(=��)�$9���^1�n�c�u�����"��b5��o6����lHC^Ml��¬���e�:fk��k�
5���ښ��zU�gI�ڼ�	Ap���� 8C�R���7��
1�s��l	5eY]t�� h�K&�5�y�;M���oC��ʳ�k(?�\��^��B��0����4J�2F~8�;q�i�8��'�P.�y�����}��A�/��MP�/��6ާL�$0KHd�����Sh/sW���lO=��픓8w�S)��@���������m'5W�ШU6�(��<K�B��<�q���L�{5k焥F	ɶt�*�x��'�6lUR}�i��N8���)��i�P��]�ff,�܌��Y���(x�E���G���3�?�NT��'J�(�4�0R�}����'^����L��E�O�
�ٌb���{��%[�/�D�?��N�+���f��M4�S;��!��*�#iL�,��|]���0yv0�-��w�aׅ�N4�#��A��y�N���L����L�0����I�����-4��rey��������k	�G���>�gKD"#�V��-&�9������ʬ{�g�:��a��@��W����y:� ���{A��c��55d�y��cx��2M��)�� @�<�"�n
��Z�S�"����D�P$����~�s����k[�f���/I��]h��p��
	�`�k�.���Qں��y��*�]+�n�z���������S�Vv8����쌯p�5M#��K:�(vG���~�Wh��b��$�fj>q�^�9�4���;�� ������"��^���eh.��b�Rz�~�?�Y߈��c���F�W\�m�G�A��v30�ٽ�_uS�2Ҟ�!������:�b��55�7�ק���A����Wvd�����˦ܣ�G�p{u�7+���� �S3�j�/��H�/����hTĐkt���3�Ɏ�P���	�gɯغ�$�F�C�Z��tA�8�Ԣ��΃�����ք�z:�tR��X��Q��!D������B��S���^(9��˒���ES{�R��B�l�D����/�b�O�`���|65}{�g�5h� �t�P�.2�:!, �P����W�,4)f�0�SV�b�3��)���\M����-�"if�*#�^�æ�tqy3�xC�Ӳ�^sh���x��C�1w��7�R�)f>�K�"b(���/�?��#k$���F[їϣ�6c{Q��r���v��(l�\�DL�|��x��U��Ж��|���ƚ��t�1mlx�b�+�����g�ea�	Jr�ӷߤ6t��r�TNb|�r�@M�оV�o #v#�o�գ2U<Ļ-��؋�#��$�\�����C��g���� ��{!�dv����6���3���ND'D!��Y6l��(މ`��9q��<�~�$���@/j?�����'ԇ�P���(VOmX�nO&��G��}0_����չ�tв)���[`���냮�/�E�Ú��R˚�<�'���E�T�g4���h����F~�[���0��%p7�Q9ک�H4I�lm_EC�8��k/�u4>�ڻ�v�D<�Ό���;C]��>lC#y�]/3���[FK�a�m{�J2�-�Ryg��u\�V??��8�E-�%�w�ZKæDd�}{�Ɓ��a���Y.���+H�� ^�߅���EV�B!Qg��;�7gYv �HqP�q+c�
��6��VD{O E���S$������	�6q���a��05�-<�9�4��o-ͤ�h�k(�[.ݠt0>Ʀ@ϋ�L,
�I+�믚�-b��?-�9�B$�Yף���´����t��ސt�xD�m�r+��0��ӆ��x���3!�cO?��l >J �BKڌO�Q�r�z�(H���,��Q�ô+yֈ�$��NM��ߙ$.{�Od/T�k&Z�]��ԣ�1��I������}�:�ո"WU�.͠���,�9��~� ,��a�b t	�f�gY{��/6J��ač;,�++�Uݞs^��xmd�2���Piz�|��9��6�OU�Lq8�5$��م�Y9��,I�e�.�)�{���L�R��.k���l�xuN���6媩 ��1���T�+4?pBV��C��
N�N�f����,P��b�N��3/��v�}�1l��߲��r��U�}
�@C��0�w�+;�)f���s5cz�k���
 6(���|���mC��M��F����ܺ���6#�7#_$��eA����0�Ȩ?�L�v;�����V�t�8�Ox�n�N��8��L�	�p ���v�^��V`�ޕ��D9Ecp@xܩob��k${~�3��\wB�T+z�Ζ�HE^��;�U�&��)Ӈe��.b����81g�"%��Wb�N��!���i���Atj�L]��X�GB���Z���g�/�#	�2 ��I�/V,�*;B��1��q��2�U��ho37��K��M�
�W����.:ހa@��_p�|���~�D�F�a��=zǭ���p��H̉:UVST3U�&�A�f��߹�kaV7��&�>�v���~�"+笧�h���ʴ��꼪��%����c��D���;�oZGL9����\�`�;^���%��'"�rr�+C$��%����Ѯ ����]]�J����Uv�V�B������I������mч$���#&+�h� SV=cP�S	Pf���T;)�J*��mg���eX~ƻ�Is�k5���+���Iړ��̂���[Q�(�Բ>_]u9l�8�4D&%m>&48�"X^98�I�|ǲM�3���kB��n]k��yu���m#K�|�p��<C
�f協(�{�w�6@H�/:��G~	l�M��]�R_�Ý;��a��W��mq���M�H�
K���.�F�C�Ίe�#���7���~R�Þ�\��!�u�eX�T{��?��O8�
x��� R���
�ڌn���;lS���8S���&G���韩���3-B��Cؓ�M�X�'-��A�8�h�2�ǻ�y���r~�E>��r���:x[�1u~ �S9Lێ�t��V�l�>�V�P�
�?�QƯ��m~]Ӱ��<鎅K��A�J2�~H��s�A�����#'���q^?c��KH����aOYfA���9�~S�`�@���x͉2�?=ڃ}�ƛd�&�ϧ�w�s���r���}�������v�]�MÍ�'Uc�	�ny�F�ZOb _�0��)�\��ە.�?��_A��^e얂�}e��=�*\��^��{�� 2a���ಘ�`����\���'�q��p�3~J��s�+W���t�>�����l��7����?![���a��r_8� $"��I��������~hl&e��_�{���#��ܩ���ѕ��c���.a�h!�� ��7�>��7�u8v��St����ː1��E�C���yv#�@e�k�CqUGEH!�0���j��� Hv6I�o�A�m�t�䛼��<y	�b�����~�i����7��)?R�-�	�^λ��m��һ�����m#Hl6���m�c������������U�J�=���Z.,q��w_18}l!�_z-�m�}�H��?�MR{t�mC�(�̝c�N&�' T��S�R9�'h�٫0@K㓼��Ҙ�
��xp�o[���/EL{w�۬F>����}�3)�Owc�7늼�+��e3ۀt���#�V��f����bA���Y������L�\bjtύ ���W���	On��A��׆¼T����Y�;S.��I��ל��a�����!�ǚ���� !�(�fy�S(��X�$��m��ߒ,�
�⭥3�����ރ��k�\_|k\� &�=��H�-Ei��}1֓H�|��ef��kkLQ�P��ٶ<1�μ��h����B�_)��A��U�"u��r��u� a���E��?!g S� B�n2��u�m�,�^PP�p`>��*�q�^#�@�A��u��RH5��.��u;m���c����\6by��qe�W��u�Cs���Q��tK���������=Y��$�d���Ow{�޺�����h^�ҕ�vࠨt��y��{�,k��ZR{��1�S��K��
�U��D�G�r��
��摧��)��"���0I��x!P�;v+�x�PZ�-^����^=4��N:�i�q�ߜ#������C[�,�>�~wV�C��46�9���m�e�d�t0��E�δH����Y�����N��I.�~(�>���b)�}���K�����U����!	�u^e�&�S+��Lܣ���f��ڎ)X�$� �j`P(����X�鳓�i�1�ݵPf��+I�֐��1J��^/b8�سT�`�A��!���X������XҎ6��<3�	'���I�=�&��+i��b���<��]I��ۘ+B�1��9��G���L����z�����RԈI$��� ���%�Sd�C��S 9a�|���d^�����	\}�IlX����К�+G���j���!
�G���,0�tS��JM8,ԍ�w<���1�z�ܳ�q�d'P��bo
U-s�S�V:td��P��2�4,��n�⮍�g3Xb<U��K
���C��+^(EK�/6�!����lgu.n��kT��/�yY�L�$��ֲ.]��*����aT��wQ̦�E�#&��2X�'��]˦8.��O+���.�"���r�ے��->�8\���N_.Ng�U1?d�����vKՈ��8��u5�2�dG��/)�y�;D�l�`���� [|�!0�E�ϯNSrX��9\�%	�G�
�'șчx�o�ѤRذ��|E����pv�w~���2f��vj�v��驲��+���X��th����Ճ���D���V~��0��M~`��eF���XT���ϴ|�������fBTgzԁ��u�<�3x��$�g=��~Ɏ��w"��3U�Ɛ�-���!����fe�>�I�W�P`>&�-��K�Yg�����(��J-��~�P6G �������60j�54�O�~�FT��9N~E�3�/��t�D�b0D\t]��ZdM�y�;�v.H���n�B��Ե8���VaS:wO,���c�&u-�]��W�O�Q9XY�=��Ilw�c���پ�m~K݉� �<�X;�����IQ�@��_������{�7k��Pa�=�#�����Җ�'��R�j��Z��)�}W��' Ս���;��*��5K`2+�pS�bq)Ŋ�S$��zO�{
��nd��
;�AK�-��3�A
�m�Z�5ch;8��⒩��=�?�ݦ�}*�$��X�FCo~���vG�J��~�ظ2������ql��Eb��K��Ÿ`i �K��(m�Ďȵ=6��fI��҃~Z0�mS��i��[���=Y�	��Z�������K�(�G���1:�!�{���I'����;M��[�)n�7��r�J��=��(�M������j�׼_�st����r��S�{�م��
�&�w+W�맅XΌĨ!9��R��ɭg�˘���N>g̩�V��V*/�X�_��%ګ(�6�<}��s�nnEu�?�3��(��&�pK��n~�#Ћ	�i�� Q\x�@��(���x�7�o��y�2e,i�z��XW�vk��E�ڌc.p��3�R�sZ�׭?��aķ>�$�OC�őx)7AW����>7wA���]5��Թ�����>���hP�"��⾇:�J��`2�n���� L��s���V9R��j��(Ri�.�tI 0��Ru�0��O���C6�2�1O~8{0�6V�G�}i\$LVH�Y��yFBr�$ r�ƿ���ުAJS>�;�<�F�E/���{!"A�4��*�Ԟ����N�*�D3�߃?�T�6`�տ�J�Rl��:�����L�<T�Fwg��5m�cm�A�υ̩5e�g��)����
:��A�k��Z�#�!���p{�nx��I�ܞʂ짗Ӻ�Ѭ������6���Z1<h(���$���b���l� ��t�S����'�X�nD%[�S�`�+��k��-Yi�+�[`��$��T�ڎ��y�ĩ�]+�%,)Ia�8ȕԑ�K�������YBzG�4z��:pǉ)���d�T�<UtDւ�����\H��Ϭ� ь�\���e�4cvGBE���W�)NM�]y�����ڛ ���Ʌܽ��~���.���f���.���1�v=���N��^-T�t!��0�{s����E���]E���f��A���G�:}qf.���kfo�v�c	sv�c�ܟ�3ir�nV�،8Z�`�T�.���F�=Q�S*�"�T����Rx-��\����RnS]��W�N
��L[�w=0�V��/A���t������{������j��:��i���uZ�x�=8@��쮌�w�#��N��c�c�Vm����A�#$�㺚?� ��ؗ�oԲ+�6B�~z�m�r��EL˱�6�ʕ���b*�띐�A�2�����K�z$N��
�F���za���Ix��{�bZ�)w���A�2��!IO҉��5��@��0Z���޷#[�u�A{ �MV���[�߅�546<�c�9+�=�;�Evb�bF"��+�e.�"��v�S�j.�~`�{��xL��� �"�t&_�O�(���'�w�&���4D����L�󨁟_C��(���z�J����90���_�� d��wS#Mp���k�SB�5P�IPMq{Ʋ�#�t��puB�*,w�6��2�Ç�cǔ��q͟$�$_V[r�="�ԟp�;��P��-f��u6�Z�R�Ǔ��!�X���r����x%p��j�P6t�OI뢑� �}������):�S�`OhS�;����BȻ��i�#��*��q��c�}�Rm
�����,:�{�ܶ���Tx�^�yr����p�_��D�ʎM�PB��G?>I�����z�c��ɢ���#����z?�����R�r���F��ӔX$��C�%�'��P$�YwX�;[nY(��R{�kE��b� �L�)�״�����VQz�vB��p{O�Tp9n�OTuZ5,��2��p%����}А; 4���m���I�Qq����s��LJ�eD�ʹHX?�U�]�IԖaϨ��q��}�9I��'j��(�~�gq������~����of�3�.���%�KL�x��؋����0�~��	
)�^�����E?b�Ԣ�X�+��!V~�Gf�6<#I`@�1\�M�P��K`����sʀ�0hSn�B���b����.��m�X=PL���=7DϮI˫�]��BɬO��adx�
��z��.��IM�+��.��D�q�I���T�*�MnBGXOhEꜛ�Ռ4��ƻ����������Ey��{/�V�y��n���7�ys�����#+B��V@���	{
w(����?����l=���2�AZ�Hrf�l�c3#_��/X?���b����Bn�J�a���	?^�l���dݛ�F�DQK��E�U%���b�9Ҭ��R07������p�.�SQJ}�N�������hZ൹�@wZ��j&h�����e�����V9�G*=�ε��`5+vsܬ���>�N�`y~P���>�p����SU����hnMcu�}5��;[F��S�}Eq���r�<�[�'��|5ƒ�߷4�c����$gL����^��g����0�Vk���l8Y���a�||�l���h��~�ʰ/�ƕ6,�P���P�G�˂
F�y9?kʢ7-28��=k�{�R�U����<�j���SG�#�x����7��ƿa����*����\�6\���2�dJ֊z�E�(�c�S�m&����k/�._�Bh��K~W�g��+�$��ϴ{����Vy�M`!��y�.�)�S��U�vl��>�Lv�7l�O��7o������KV"k X5���"�����W>}n�����u�� 
�-Uc#����mH��K�r�<�f'4��`۰�mJtx2!9�rA���
���J@OB���Hyu�]����|3���/�`/ZO&����\�$�O��������#*	���VoV+�d���v�s;�=4��m����Ϳ3;���7C��B���
U�G������;쇘� �Q�S��׿�>wܐ���E;�ȼGӁ��U1��cQ9ח]��f��Pƅ���0QS��똵�ܿ*��!MT��/�� ��?��Pr1l_�$�o��N��Tjl�}�������T% +[��֒�>é3[�؂F�C$��X���Ȟ�#�Ř�:_g��P��e���"�?����,nJ�Q�r�₃�t�^͚��N=A���lf�=X+@�T5�WMRO��@(�8� -Dň��PNpV	�p/�����Y�B�*�YBC	��V�x��iP(Z4��r��w׾�ҋ�����tӘ2#�$�id�?����}�@��g�ƻQ���d�݅%�RC�Ҷ���e�rX������d�n(�����&�N����Ɠ�`U����
�]�+m>	�����N���i<�����  hc*z���p��6�Y8KK�D.�m �����jҺ	�������|ȇ�v4�J��<�u�m�)Lt�-�*L�Q�e����3��B@uk�B�+��ԂIa���ޫ��	td�]�ܴڲ�+��}0��@�-v����Cܢ�������e�wZ1v�E��	MWR��H�;�����fG��(�qZ�5C��tQWŜ���o�0�_{�i�> ���'�?U0��=�I�����d��+��] �����W���^dm����`b�G*k��+y��K^_DÓ�{A>��E0@��bL����t�Ox7`�S������X
LS�yC��ڂFdx�HŽ�5�e�=��F1\��.��x����W��Xs�fy����M�`����t�My�B�"�_���H����eA"�>	�x.����Ha��\y�P�Ϋk���0;��ݢ�a�5>�TY,����"���ޱ>����_S��>v� @���O�Ůa����k_Z�6�T����}z�<LEi?jVb�pK�F����%�WiDӟ �`�$jD�����u��.��^�;�@i�ol�r�e�U��
F�ք.E�X�kS���?�|~��r�ܫG�Y����Y���.�X��Hd��iT�����p��J�����vN���q��e{~K��Q��8�w��w�K5Q`�X� 	�ۍC:'o2^����/ױ����G|p�q�n������苽ф<�lC�J�g<[��
vQ�'	�Kv�E;3ݞ�b$�/�����r�P&jh�%Xm���L�n�6�+��r�H��Ge<�1@߫W�_<���B4#������'�l�,KWFy��}�ץ+n�n-㉔�s䇽��(~��K�1�-j��h�)Or� ��EJ�^m:��f�R�����YҪw��gqx��9F�<j�R:v.�(�R���6�v��-�X�j*a�9�k��G���q3-4�6T���F����Ѳx�:a��Y\&�l�m��:�/�,ѭ~4�У�ӿ�ё�D�A�,Srɤ?�+P��u�7�i�{�v{����h9�IEf�֨�n�4�yp���J4�+<k�p�f�	�tw�|~}NQ:|���MjNNΈH-��~#�.���<&wG;�c**^�J|���^t��RAuzw�-���'�i�[�	V7qyI�����'ke�� X�B�m����}'}Lk��*��y<e ���! ?tXj�7Rp�����X���z��i?�:�/�()�o�6���2TP��^ ���Pb`������*�{_�ӸB���wk:jX�M }���u��#h��SU�/�H���h��1���#@�u�?m�O����-S�2/e��7#��*e�[D�1���r.����N�j�+�tL���s�H�I8B�ٜ��ډH��Э�2������<sn�"�T�\��G���J"3�M�𯅆I�����G}�=yo��t��V��~��mK�ꖯ�[3G��^P�E���j���
-��h����04e"�{t�,?��Ҿ���������*e�4��M�K���������
a��煑�P4��h���S�,�o��X�U�3F��D���7j�L��.���%N�}Hx��RԖ������;�;�$�J�Q��?G�嫪��s;�S�RA��������
��Ai�#�6B�6����xvDv��~(+,���0Tꯌ�
Z\�e�|q���7O�<�Y��@��i~:v5�ٜ��쵫W��S|�f�(�{K�S�-�~���u�7i�ͼ`���BiZt!<b�jx}G��S~Z6����^3��ߵ����^v�����@ҫ����0��"!����v�=�958.ku���ܤK�y��ʿ�rn��,�MGK�7�O�PC:�@��)ᛵhFԬ�|kD�m)�O懜V�xJ����th���g��lac)|��3�����?��#|�Y��9��'2/Bfm�ʍ
}�#�^�DX�����wCS�XN�,D���_0;W�
�O��� ��`��
d�U�4Ur������*��G�3Rh����tު_�u�ctG�J�Z'���W%���?��@��� � �A�?y��E2Aڏ�(�s�/N \�A<a'��6��҈S) �NM�ma��b��;��1����C�g�n@�WI}�Ti�\F�؝S\Q�W��]�"�Ov��_߳�5s�uPD�=���dR������o���ݺ��*$�^���Z��S4G&�!sF�D���s6��f2�_�BM�2�{��4���@��Z@�U�G�`r�5���-���C��3+eS\ n�.�I�����^z���&�O�ʟ�L
=w�L�+��]ٓ���Aڕ9+%�l��"�7\��a{9���� ��J�E�A�4��Щ����ŵ��ы@���,���;�y�\�C��[R��Xn�Wу{������K�x�0�m�O�J���F�k���փy&�C�Ĵyja�5��'����)b,�B��L-�f�x�x#�xa�+�E�зk���ꋫ�wS�aX6��R���BE�p��g�o��W�W"oK-ї8�jt���%Q�&`F/v���2;����нM@�']���ٶ�E��4w�ɐ�@�E���F���m��ے-"�`R`6q�4�ZBh��ǥD{0�"k�i����v�����D�ڥ�8�Ԉj�D��ܑ�x��|�u]���؟��h�S�%��5��jqB{QZ�1�W��h��l8r��;6����X����֯���`��?��8�k܄��g_H����i4���#Ѝ
�)�� x�P��E&�/����*8���ޗ4�����O����F_����'z�A����!�?�Z˃��c��<���b2�^��m	+JK�ө�Ȅ[WC󪑶�*�i�m��d�8��W_�ʧ�GQ;�5���E�ā��c?�G�H3�v��F)��8Q}�#Q�%��Sj��!D{�Vn�p�v��%F���揔�9R�\�H��$���4���E��m��Q�od�������X�Jӆ5W/~��ٕ�o�3,��bd�?lF	�$J���;g���F9ʫ\�#��D�8`�l�:�i�Ng��qׁ��J�s+/��X����b#��,�-�Ċ*R7���E_NVD�y���m%/�/#�;����%x�N\��+Y�g2�r�1���
f~��Z��ֈ��k�z�M�΂�@ϻ�9R�ςW����_|j�Bζ�yvJs�?�:�~�Ui��4�mՍon�)I�]4DP�t�+m�&q]���D�{ʔw�~7��'-�y8`���H�0���r.0e��q%5�psFr���ȓ7�dv����P�	�M�;��n�[U�.�ZI�]"�RZ-���z���e�JUy�l(D��C,����j�\��j� �11$�s�� ��AZrئ���|,5�5�7�AYv��/D��!�X�����-�L:y�?�ٗLHm���b<I;V+��O���ɶ���~��i������0Eu,��{�۳�\�5���~ݱfV�7��{�������|5��Fn��FuAJy���攡6���0�7�A�c:(�u�*� 6
q0���]�t0�JW�o(���s�_
�IBL����PrR�h�V�ZbGj�a�~ng_�:��MÊST\�[ox��}��s���]ٙ+�<ejg���?BJ��Yn���.���ca
������+��É� ��B|+��vc��5M��M4�,�) �(��y�Hޫ"O��.UV�����yX�R�(�y�c��1���l���(�&V����˔�"g�n�JN|�3򣽱�k���aϛc�F�U�Voy�h|.�+#=��U� ��GTdE�u��= ���+ݑ쥪<8��+�ŝT�r1X�	q�X�,0��=R�x�c?\�@�$0d<��Y�5�kP���7]�\���5@�a�TP�'-5Ss��MS5w97CXD�P�'�qK�qOJ��6�,�o�����0��5�}�Vh���n���Q���ͦ�"x`�XeS��7����O@IB�Sq�6�k�kmJ�tF���;
�N��F���95'l3 B��r&�UI�}��~�ԥ,�(g�\e��nR_�<�����w{D�$F��sCX+����u5��%��/��?�"M�Z�x���<=	�:�

�I��	��f� �މ���5��m�Q���g���C�f�4�{������u&��BJ��=>�ϱ���c�򉹊7�Ć��c�Sg�1����߈)�+��&2��a���Xt�<�F�y )�*��1��P�CQ��ubc��f�&����gChԝ���A�)4��U�-a�����z���EՉ���\��e:�!l� ay�/���
���[��!�p���\z�����0���,��_�|�f���B��E1��$X���Q���g��>������.!Z�:���%l��j��qjgZ���jT�֧d.�� ��7��i�|J�v�\�/*+u�.fo�q��o�����V��D�(���Io^�Ǝ=���_Ǹ���3!Zs�l��p���[b�vB��ۆ�Q��- �S�r�������^�t+�����~�������W)���<HD���p-�APH 9��&%]ߙY�i�M]b=�'o&�ڀy�R^SJ��,��eX��q�5��2F���*n&fwL@�w���I�T���h}��SI/�ڱk���{����?XU��k~;F���Zļ.�Q�E^�[��˱�������;��.��g�l(>�I��g��Q�X�80��,�cZ���}W#��b�S4k�Þc�{H�Z�㩋S����&����~��N=���N��U��Kz0Yڝ(A�z��3�q�^�������P@rg�]*��h�.}�[Į*�������j����|?��"]�V{B����0���!�t�.��|(̵�g�.����T2�'9fד�Z�[��"P9�� ��A��g��At/Q��>�~ӼX�-R�W���qԏ�̚�V�{��%I��l��<8Zv����G�UgccDMc�L,E�:O�(>��������>�߂�!k����)�/B�����(�K*|�7��0Li嬊�)ơK�8f���X�t糜zd QЫ��%! �H�ɷ���~��^*,�dJ:�˗� vBV��~xY���� i*�7.�B�A�hb0cL��	��/���b�Hk��y�&pdb�e0|�Ҏ�AN%�z���q{��=_g�+^wS�	�<c<�j���%��0A���~	�>�[��	[j�۩���^Ѝ8�4C�`�Plq�e#-Kf��x�H��h�T�����k'k_�Λo�h�K����,23��'�$2a�͇*�{9�:r�ru�4���>����0�ɰhD��P9�������I�
YVR��i��nI)T���z�E��U�cH�Yt�6��H�ۯ�� w��M E��[��1N�D�
(%̎z-����I{	�VL�i�v��d�c�O�N�F^#m�~���bE��I�C?X�=HZ���"��{� �ܟBv2�c�^��H�Y	��e��~$D�a%o�-��(���?��%�9�q���|z�(tƱ����#0l��S[�����I�efP���A������,&]��?ŁU`dt*7�p
;�b��-�)lV���Y|a5��Ȱ|CR�~ndeTXT�]P�R�3r��Y8ڶ0�6�j<A��~*�`24$�H9K���ewp�kG�\|Rjz�M��Q�(o���������T�Uc�	�`=����%QtH�0wBQ@�H����s0�p�Wi_�:�Ӂ�tR����.kv� 9���A��w7[��!4�K��<~/V�����|�����-R��j�@�\ �����D]�����8������D��,2 ���u�ٯ�k�iO2U�١rգ�"r5,�[D8-II���UZ�ǵ�=�Z(���&���9���wo��Jɗl�wԞy|Q�#��u��GR2_��f�,����\m���{-�w�3�^cb�
�F3��o���,L����S�p�<�a��Ij�����0?��&�JW��8<b�_��!���E�+�'l��G4XM�]z�ϼ����!�ʣ��I;�ɔ4�t�\T:�&���mGr�lF,�B�r�+�isO������\�4��a(޳�VN�%K�J���0��j�B�����/x�SȷR>)+�E�<�c %	7 �v��t�m�u�$`��k���DȊ�N�Z*[]Zi����nS�n����n��Yݥ�2�����G[V�_����^.���)g���s$��LͯAz�i�N��4��/�-��gVQ�����;e�K�?��V�B���@Z���J�nK(в�ye�V��H&PV
K�<n���o�
yy5�m"o�^(�q�-z�[K�	��G���ޢCV��hB�s|��z�����#lz�gS�9���.�0R�jK)Z�N7��@3o��2(�����>��Z����C0H.���q_U�I/�B��>à�X�9��������G���/c ���[C�uj�&>m��mg��� �s��%�}�$�nK#.��{ T<�	գ鐪&l���:~%�Y���>x���{���9�%Y���*���)�ɿm���H �w�|A	�>�R��i���*~��x��P�	ta���&�4��1�J.'��;y/U��7%�����vѕA'�Pw{��I�� k.�@W ���~��&�pK����Pa�2�%�G�1FƁݴ$ǡ�R�!>�qg�?P�v�o+�Y0�_)��u%'p�v�%/��媋MV��c�[����иʘ=�I��ӶS��ſܮ p���w+�WO x��LT�>�?��Z-*��4D�ϑv���!	Kh�9{�u��i��<��7�*����s�j��{j�b�"�:�>i��4�-�\�C�|�j�Gi��>\�V��"���~.�?�$fh��EP��Q��s�z�5�t��/�9k*0k�r}�j{��;i�-i(4h蜳���Ie�2�{5Ƿ3=;��ow�����c V�Y�=�/��X?X{UXV4@��T��x�@W��#����ZKiD6��)�}���;��{��yVI)��n�E�K��R�r|g�w$is��@�>�`ģ?���Lv� 2�F���AVcCx�3 ��I����@�Aw�F���P�j���[H�>��	:	��C���� �S��A6'���H���1����M
���K �e��{<���g�$3uT��4&wȈ�A
:�#�]L?m�0�m�W���?�����H����F���g��il�k3�겵B�OH!V7��J���qO1�9�sε������o���_�ֶis(�v��)x���ݷ-oS����w<OC��T��KU���NY�S@�t�u֞���� ~&u�
&��:����ŇGc��RL� B9xc��~��%
1"�<+ZD`��+.>5p������m8:�"p���Հ�r]�"$0*�y=�
 ��vq��e!��\�>�?;*�jRek�@d`|�#����&�R��Y��#(xS�lA��v�9*����N�*R��ob�*�#��3wq��G�;w��V�n�a�q`��-��^O�n�1��J}�&FN�g�����x;�eai����X@��]�Yt,z�mQdS�٤�l�+T�5I�s�]��2��ΐU���1��w��+,�(k�4Hw��s��1tp��6�y6*	i���M�,@�7��#��}�\n%8O�y���_����R�ct��m-�j��c�%mb��{4�q(� ��ʬ�� q7d��H�"S�ysA�uM�t��[W��ݨ[���X��
!�͢��vҎg����������Н���^&��/�c�]��HU2QV�1z��zU�@���֝;�С��o��D=Ԗtp�����0�;��S�؁ Hlxaq��%�ǠD}�ɚD]��;����)�W�	Q`�e3���	j�4a<����VlS�3'��pH�n��3}�<U8�w�IT���Zm��,��S�N�i\/%7�� X�֜m�e�&���#��a.M�L��V��J���~�~�����B��h�s#g�k0����5�BnXz�ؔsɽ�?E�ś��ua�p~d@���|����)>���.�� J���O��Krs���}���'�e�yw^�0隦SΑ���b�ro�'ZRZ$l)�n�r4�0Ǭ����4��j�2�7ӕ7�`1�]7�� Q��Rܷձ�-M-�IDe�*��74�xŸ��\{O��rO!��Qg40�5�׎��}*�+G�S���YQr�Kx����ǐc���Â���fib�I�],Y�rI���[�Q�/�c�j]YG)=4�Z7�o}f�J���rɨ�ze�!��O��43�ɡ�l��B(�d"S9�6�I�.���ˁ���̹��T=���T�����H�R[=G��7��%���M4�D��s�����XD�מ�QE��a:ԟ|&�WҔ-�[��$��>^L��Q�뎅�d�1�o.d>��f�^` q'�c=~y�޵�Y#kJ�$�Е#{}"o��\~�Z,������u'���*	�Ct��e����t�(]>Ðz�?��u���2h$���y�9F�Do�I( s�P�BO_ɵ[Ei\֡*�zi�L츣��j2��P�x���׬�ɓ����Tn�fk�e���I4��F���S��#�8p/x��W�^����|Ӎ)��ܭ�L�A}TH�z6g���P��_�ޮ�E�?	Z�Z{�/���.k:���/_�����ne������`I��|ބ	���6,�˕�O.����k��+.}b�[�Z� w�8�v5��WgDu&��@]�6h�׺,���vG�`.����ҲfZ�P+瑥��e�6"T>d�}��ԫ)MH�x�҆�wmC�ܿS7��������)��^���hP�gG}��N��U����\u`%���������w��Ʋw��e�ճ�O�������?o�8��;��v 5�|*�X���@*��7n4���B��aςsm�H�|R	Q�s�J����/����j�~��s�0/k�z�`�Xs�B�v�Z�:��?.�[��a=�>�Xi��|w؝	f���6b4��u�Zn��6S�B(�� �6���������۸����)��2����#F.�?�$.�$֙�=T{a׷�74.�Z	d<g��O�N<�JҺv�� �6�	�]��?x(N|MKw����ϸ3rͷ��Lɓi�fœP���y���j����AȂ����E0��#{�IW���Ԑ��x�+@ނ�
:��Bf���:K\���aW�������/ΜB��< ��v�
5��qq�����D�m/7�W�6 N@^����# �fg|e4<(֠�k{�e��ͺ�z�\&Yv-k@�U,��$nw�f2��*�@f�Ј��Įj����w_��dY�?�+�����c@�UV
#v�q>�}/Ƽ!{2�,{���HV�#��@x9����Z.o$?f��5��C��I+7ލޖ�B���E������>o� .D�ldk�pQUT�!*K��U�'m	\0A����5�F��a����3Y�1����g��u^�h[�|������ު�h3��wyp���S�I�F	 ��G�^.�R��򚟷����19�B,P��9�P�ͥA�c�f�d�C�lxg��5��kփ���M6�F�M����pE�����O�q3���S�Zs,�~)���LY<��+ =1��E\[���<��$�˓���	@�l>��2"Y��ǘ���Y���Q+gY �v�N�]��t�@�4��iy�M��Z���p��qV�mp�g	��6�d*<
���or�ʴ
P~?�H!-�QM1:�lLpq��T�q˿��f:�l+.�>
�M��@B�艺�>OW��=4T� kk�fl�6w�nR���ѯѢK�I��2QA��h���OaȆ����7LA�A8d)�qp�Bdd����b?`�S�&&B�Qn_�d����Q��g
y�������=dc(�ͱ#�g �n����w"�-���f�3?r�r#�ǈ��c��=���:a�.�~�Y�D�֝�:!��5��튕���R�z<��a����^5�O�g�Tm��d�̤��O��%$/DPn��-v���������Tܖ��T$Z��瘗r
��D��5��O����\����*|N�zxG�'A���x�]��X�Oo&In�I-�D�g^�p3��ֆ?N6������7�����'�y#ǘ'�gF�A�R�Ħ�j���D�4L5�p�3��"��;f��Q���ɜ�)X�'������%�F6g���Zm�,���D;�Vd�YQ]t�1u�:�r��=4x���q�=���5����ΡIA����j�A��"~L��IAk�Q$UA�3���__�](%;�m�Mp�s�	��a5Θ��HEwӸ7�'R">�.������Z�;��	���~��]�Â�S���t�E�,,���4�T�ʆ=K�I���/ohRp����C$~R��5�=�z,����P��Y���d���� ��˕v�x9+5����gN��n�'s���Xj��U�'��Y\m�?��1�H���ʛ�E�@fo����[EQ��myG��
��g̼o�<�N�=[�[��3�D�!Ba�1N`ŗ�^��9���:����FFu�hSv?�4�d#49����������h`�b�����ށs���]�o�>��`"j�!�O�S���0��t�DqF�K������T����7�s�60A Ufm�v�?N��엋���M�M� '�Bm-&�3U#$F���av΍�7�I�̕������69��X���H���M�hA��4�}�Uĸ�8Z����#x���>+n�NO�	$Ơ��L�)��@�ZT��`��ɑ�x�>a\J�����J��-^"�����w<	�:4���D����3n�L)�h�K�K����_�ydڌI�+���)�˔Kߠ[!Ei�`a2w��^k��H�Xtqֽ��Φ}�EFk��|�f�T��5�$����AmE�c�	%��e*]e,���T��Ou5�T�2�	� ��l?(�4/��I4��D�ob�3A��.
�������\��������x娨z|������\:�ᐸd���,��⇥��?�zS�܀������|J�����q�65؋�р �vu���H<�^�	n���?޾A���?�c�8Q��K$	FeH��.�}*b��0R��*�!���u��E*P)BG�l�����D�dN�Bj�b�\�8`f�0�Yc�~�`�s?�h��L���{��L��EH9u/�����nٸ�?�wbbMQ*�?��GzD$�ŵ���)Έ���d���:zF
�,.)v��Bg�겝M��� �8BÍ��X���g�}����T���:"��[ ���A�d����'K�vG��o,�0�����ߛ{!F�sJ�'���iZ�ҠC�V��H�d?���sޚ�B���<���r՟���ܙ� ��,���Ap�w����3]����ģ8H�G��� ��r�x��zZ�����s��-U���M�*i���=��(�p"4��)^|1��Z��st�q��2g���֞'�$- _6���*#v7Q��~�n�O�[����Qv�Cs��2QK�h�mFmӮ���б��!L�^��&�DhiZ,
m�rs֭�y�'ѳ�vr�s���p%���ԓy���=�f4.�4�g�*}�z�"�4����<o+���Q�#HI�����|'� ��ɸJ�%V�EU+���)>��JÌ���M���W_��mEJ���F��0�i�:{D�G_�6���Xyҙא)���L��̟,�7=�=b�S��=)���E��4�~�-<Dz=�� 1��X���p�|#.w�@��D���q��� ����I�?�m"�u]�����e@k����)�H�0��1���ʞ������kw�P1E��4jl'�LJ��4�Q� (3B�M:�R��R��M	�����vY-#��f�an�^�8��-��l�d�sy'���R"�a���ׄZ�0�,�J�î�H�Ĵ��o�<̑m(o �[�Zv�u�SB蟠����N�;��΂�f�ژ-�L��r�&owa�4���a�ɟ��i}l(���:�L-�rr�J�L�v&Ԇ���4c$��:A�*�66`�Ö����h�8��b�R��	����St i��IwgB���f.������Q��4u7|"�|n�|�iS��|�c=kh�ȧ���H�q�\�O;{)f��qa0.�����6��2=�t�����>��ʈ%�6��>��G�P��q�s�/��.ct,�
��I��<.�H����=xp!��8) ��Ű��(ߘ{Z� ��v�	㟟^�ܡ�r�lQ���K.{QS Jn� ���䡞�M'w����.��E���~C'n���Ir<�}�0�n�����d?�f҈�^��4ČmJ�&3��7~}˝<"�6���Zb�v�+���7��"P���d*��e>�6��H�;U���]槩UJ�z֝�h�U�_'a���E}�"�m^��
��+N^M��`���?E��:�H1�<����9:L��Jz���~L�7�)9U&<�娓�i���)hc���CQt+�a����K�3#�W'�`d[q]���GP�����V�3���,���h"��2�j��_$r
xRL�Qc�v�dK�kx��0�;�x)��:x��S#2�i��`;�$(u���?I��W��cB�����#�s��-�׉���.+2���/u�w�Q4��2��p��� �����>Fk���3�k��ȣ��xR��5(#%>-"XgS-�����>�<��]@ʼX����)����>j!f��\Ъ��m�j$�쨀]�8	�P;�F���T��{_/���8	�?�ޏܖ%Bcu��=kz֤�[�
�/�O�\���t�4�'&���Jc�GOnނk���Ʊ\�^I��\���D]�*�*��ۃ�J�3<P�XY�,�%�!Nb�V
��~���ͦw��&�R����9X�?�*��P�����S�.���#䫋�5�ؘ�F%ڂ%��ؽ�x���~f퍅4�Y�k�N�)�a�!k�g:Ii�Gcf+���1������@�X�껴�j7�G����CQ���}���j[ֺ%˰�B&�dt(JE�����D�X����>�k��ŀ�C���M[���nz�Nߢ5��'��Ùt&MK��^®FL�&yu��p��\,#��i9+ad������m�D����p�]���F�>�Z����CB�F�*�`��R��|��ճ	��#��r3K�l�B��PL�X/!nϝd?f���I�c��'d����>���#t��h>ðչ�"��D�v����ы���s�w㰲@-=5s� ��_�QҲ��T�� z�^�2���rD�|�#�A��\Fȭz�5�X�'|RCR��m� -()�c� GF�Ĳ �vk Z"�S-���!�j7�Qmշ�P�d~y缗�mGm�kd-�z�k��W�U�p��8	��)��#��,������Д�m���<��b3qu�׮��V�Fg)Bd1'���/��o��.׌��l^
ʔŬ��ն�6I-ֽ��%�V�N��^�JX��1c%�6q5Cy��=?��&~ky��6�9�MKeRrD����F%#�=�a10L�o�1ms�#?M٩���pd��Ğ��:���'ک|7b.�
`��)���-�Ħ(�&����6��%֞g�k���iݕ�Q�ݾu�%v>\�v�i�{�B�NB���B��*����!lta2�$�oŴ+�7;��|�-b��9��6|S]���rc7��/#L\nL�0xR��N�k��`�Ok�
�m��I2�lk��)��ċ0���dٵf� �	-E���v�&1���U��a@����׌����hٟ)�>�6��Fj�z�^.���q:���ׄ����v��;�xꑽ�R�u�W�S��b������.֩2�f6��o�r�M���Ș$����&WԬ�Gm{]Qe��o���I����cLoE��W6�|���;�c��u1	��}&{����*����E�o>2�t�x�Z�r���y��h��n���H�T8�I��	$VbR��c��2̐~�|l�ky�Q;NQwR�n�'eQGIB&�I�	M��z�_$S�'b8k
� ��c��'�!U��o�&D��/n&Q�(�d���i�z-�`)��e�x���9�Y9�<����4ʰ�I��6�#�ac���6`2Ũh1'��ߔq�����z�&��Y�n'L��#.y�Ț�+*P���m�a>���
��'-����W44bD�]����Bֲ���L1��4V��}�n��$��ϠU-l1s�ȃ$a>v�K�J�ڷŁ���60��z��w�,����! �����Y�ύ���)�G�cI�� ŕK���3K��'R���[8���^���3d-Q��͋걲���^�O��o>/FIR~�~d�-V��C9����
�*�k����gU�6�B�;�$*Q�EΛ�un^jE�~�Ϲ��0M�^���<��͓��X�G�� ���W�\����#_���U �|.�6Ш��Z&�О#����$�2 �+��O߲�0����ʴ�r�����_p��§�Nݞ[�Sh9ο��;g�{���>A�JP\,�-���S����`��<�/�>IɊXg/UO��~��y�sS�Ǽ��
���Z.�\��UM���B�>��}�s7���a�NC�|V����R����ƹoxg�v�>,�:>�j����yY�tV�~jH��g� ��^]��z
�]�c������n��L�M?=*�_%��i
-c���I�Um����G9M���֪5iK��JT��пX~Եz(��(~k NW��_�B�a�����~e�k	��*jw���z�B��U��K���`'8�&��T���8��J�kr3��*��	4�@!�C�<��e->� B�U��^��0c�i�+���Uo��tɂ�F�t����g*�Hg�^ ��{d��!����nF��o0_ܑ�D������d�=j��[{|�(?�48CB+	��_��}���`������� x;��~;3�2mҔ��f;��gJq(��W�<&$r��l�B+֯:8�U�c�,��prS}G�@�ɳ:È�\a��A��������d��5�\,/�5y��2�(�7�\�$'�o����e�J�n�l�1S��?j�����u��#�`��b�I��uE1^�~�F�7�v��WV�%dZn|_s�4�;h�Q	&�q��*�~�Q�徦W4��ʍ�Wm�Zjej��$5d^�'�.���<bsg�����-� �����ɼ��e#����%�w3���ނ�� -N%�Y��nJ��h���}9��Eg�;
�������6I���qw�
��Gh�5�
�+����mq�z�������;�:�
�W��$�t��n�f�Φ2+�K�<�i��7�{GRb��������}&�̀~�.
����0	6�\��!�)��;L���C^YNq��K�p`	ŋL6��8�-6�;$&�Eԁ�Jޱh��Mɧ'ep5�LK�B	$8���������鏹��?n��$E�k��-�����!���?�|�H�qTR�`�E�2��:��ß�(�,���C͔�7����fAR��Ӏ.�z*��]��I;�
��BW��Ʉ˸�@��c��Q#v�\�f�����DO�U�ʡ�T���{᛽]<���Q��'����ʏ� �"���ß�=?�j/����L�q���L��,0�`�u=j�F{���� ���+ �����uj�%�ޛRk�B��p�H����,��B�$M�y$=���n�,ݔ�Y�\O�;gd.7v��+#���):E�yA�l�P>Ws>?�,��CMPB�H�Ht����J�B٦|�%�z/�����:	9�m�#�(��p��� �4t��y�����ǥt��%Riu����@5
�pۼ�Nn��e�vm�NC�0��e�h���I7����[�Iy���ߛbf�)�kSJ���̮:������ʑMݢ�!�����I�j�[��~+������5@S�Q�R����]_����2"�%�q��sw+�1��:w̱�T�I���?]�%�uO��YN�?i+��t.�c8x�;����gs��E�>-� n����%k�YE��5һ��N�/�L�����?�.$���7 ����-�ѫX��'Jr�k�#oCw�Q���ؐ���A{x(X\X+�t���zW��k�#�49)XFx��H�+�����準�5��z�Gww�M�R�25'���{� y�3����p9;�-.-��_]B;Z��2����+�=��	�5Y��`�$Td=��@$+��ݫ�!��mR,7Q;��#�hw�v+�r��Y�w<?���_;�2}��d�h�7	m~��q��}�nTy�u"�$�����8j�v�)#��WF�w6�>�3?�%�g9VF
�����4xAđ�r�܌H��#
"��5^�9<d�[p/���훣O.��O��:���_�_�D=�ҫ�lɅ)n5<U�y�Pqk��vEpn�1�]u�L]L��Y�n 7�9�=�O���GM=+#��^�%���d��Ֆ�k���-63"�[�ż՟@�2��B�L@t���3P5��U�5h��I�g�>�1!��O&�'�_�տ�yOp�!_�9 E�Q�yy1��grg<�?�>�R���8�jT�0[Zy5��p�L�e[A���{�o���Gl���*Er9>�Lg��ү����m�(p����b3�f�T��{H��9����L����V�%I��e$�=�,�����
�?p�(u+�U8��\ֈ�;U fS����v����4"eSD[R�*��s��$�SYސwȦRˢǂ���	��0w Vs�' AɈ����$���g�jZmX ����r�Z�ȡ���8؂���АK=˭u��a�h�k'>�{���gIo゛|�^z�p:�,.��ۻ��H�ئ��.&B�q�FAOCG����W�5�"l9ϱ��C���lZ��u���_OxL����ϥ��D��0pR�i��6�>�OINv��{kA�*�����E�j��5�
r�+>�В�]������� &��;�7�	� � �`�� O���\}���n�p����3b������K�5Y'^���?�!1yp�~pO$������ �H:_���N����%�GE���x�s�y�eF �\��S.��M4W��n�9���^�0NY�T����4��t�T�Az���5�5���u���t�T�i��6��g'wh��'���^K�qy����5�Ĕ���K�ה�A���I墆�5��*':�Ó� )���a_X
�F���J�=p�N�R����uư���F1:`�~NOQ�i�Q�}c=sWLƗ��| B�q� ��<͟�M̏��v�ި����Q���2���'Jy@�"�}��k�x��\سy��)?�ap�#M	ꮳ��l����9(��lٱj<�(�AsѕR�^yF	ɳ�U64�Ɲ9�������܈��NS/����H�X$���H��R���?+\	#-�?ZK�k@����eΒ�����K��b�N"}�̊�m�_^;�+�?�Uz�h�o'\�w�x�7�p�����ǚ2m���V�A1ϊ�G7�-+�S��C4UT�s� �f�7yn�9d�""�����x9�-��yIi[�	z(|�/b�C��?b�^5>�>և�"9����)O�ȿ�@�:�����baO�;]R[v�l�� ���L�!Gs��$��G�[$aW��?�c�����l��v���#���2:/��=�f��2���d�u��1�<��M��,���b ��X�q��ғ�y�p�~��j<Ԍ5�@5z�~ؼܻ5�DW���:��*Zi�-/z��4� �/�*I/�n�೽����E0��U��h^B�i
�.�Z6�ȺG�a@�!0	�r��h�-�ᱳ��~�_�E|��V�yﯸߙu?� ��̺������Eam�V�ү��������MhkT7e��c~��
9�ԝ��ά�H"_hO�� �%���W��V�����p�$$�k��b�RF�XD�@6�"q	ض�~��¯P��ծ��k:�݈�Ud�zU,�hOu�q���\�f��1�G�B��pM��>_�e�er�>S��so�y`Ps�\K&U3dj��]���ߟ�QfzD�6%��p���9r3bZ����ޝ<1��2臽����f>Z��!��4�� s�1��]��H�D��!LGTi�J�X�4��p���IU,U�*���Fm�[�)�i#��I��_�*������q�l��H�͖�،�V|mq�]G��� �M�00.�l3Œ���~Uq0�_Ե�g*y/������B
�CO6�U0em�7����𥚎8Ɖܭ�Y�(��"������KO㙔i*T�ڧd>�}�Y~Fu� �@�'X�]1*�\b�d]��ȏ9(��2�c��{o)��[x�g����8�I��	O�7�S�|�8��n���n���D�]jH!i�Kp�`6�w�[Ut�U'����'�W��ˮ��b�R��MӰ�*/���x����cs�٧۝�ׄ�}�ws���w�,c��i8�@(RN5L�w"�}РG�2�d����(�+2���N$�k��
z�a���>����G�|����?�2�CZ�ZWOP�[J,��~	@O���G����Y�1�59hS����w�3�	}^1ഏ�E�V�Q��G_Ȼ#uy6��U���=&���(���+�{��i`���u�iV�����ʒ����A��Wq��@p��7��5�EX��5.%4Оq��u�Id7�*lk��vzL�M�@ѫEU$u	���8�e��nנn�To��a���������;��a!�Ӏ\�	�f@�"-�b�l�K���8H�&�7`����\��́Փ��X$��|��)뜱��hpA3j��s��1��[MvB$��H?;f���E�  e�_F��x��e=�	�8�y����d-(�yYU^Nv~�!<�7�,K�8�`������;vba����qQ ~>u��Ll�gpo%3�?��]�p�f}�;�w��?/�pMp��E��~`qt�i@�E
��W�{�2�a=|�TJ��SDX��3M'�&df*�C2Շng��
��,Z��A�Yi=YkJƠA�t�[1p��ӫ���O�s3	yS8�\&�曾���擭8���P�=�n�ך25��V� �<�vJ����Y&]��=貾� ��y��s2�l+��dc��eC�(h0�i<�dxi�.���ڭ�:�����I�֯�:�/=��'%�H��>�h��|�6�L��J�'O����q����B�즍�vm�$��G��p�Ti�ʚEH�	�����C��p���Ex)�^�|4��D�P��ήr݆�F���;��S�ç�b��PF��m�e�n�s����R�h������Sb�Ƭ6y�B���۴�ۋ4��3�~^�xU�t��G�^ :F�T�xM�G.��`_��o.z����+�Z��,�L2 �e{ġ]�-�էML�|T���P9@`�����வ[�#Ȕ [����I������=�a�����#ۆ��xΨ�V�%�aK�(��V�r/?�~m6۵%!���>j�����1� ��u)j�c�2aVt�K���\}�`b�*��zQ�؅<ʤ�6wծ I�Xy)h �M�:������iV�~u�4P�O{��=���s�"fM��?��Q9ʖi�����(>���Qӑq4e�5P�v0�ߥ�妤;d}/��Y���f��sW�����nVU�eP ���*��Mi�[�ȐY�K�=��{鬓Zt/�e]�{h�nb�d��mr�j�j����(vw�'��^��\U;�
�X���,�a֚�J��X�?�v�=���`4��e�%<�pD�O����3�#�MoWp>M׿z�^WE���H3�o{*���M?=ũ����OWƯ��6�������e����lՋ��R�v�.�dKY�?נ@3����sʫ����a���w�N��v2����5��$8��֑������,J|�>���U��Z}ʺ�6��$��hx�N(�j��%�XO@
�`�*A���4�u���=�C 0�])\����a��ݛG^:B1�a�Z�K�: �E�N��5��`#C�����9�
��(F��2ܲȠ/R�����G��k�:��כRG������X�n%Cy��Q����
[�:�i/ל��]���N�d�8m�-�y��ޤ���[z����.�*F�� :��ib"&���7�:�>���a%-�k�a����ˏ��C�l��cD�<�UY]}N�+��;��9�ʞ�[���=�0�Z��;��9�e�KF�7�s�������@��O�x�h�q��X*P:�WI��R�o�W�]�Y� ���h�đz̿��1M��T�����UIUI�)�5��I�IDWa,�}e�ZaJ��TGh���c�a]��U0?�q�(r��3��S��V���G�J+���"�1��j�T�,_p��xg�iJ@�k'πL�З[�� ��Ѳ �R[��6��(�y��D�Lt��#L
*�n�%�9�c{��r����o��)�W�_���c� ԘG�TQB�ę�����ٖp#ftQ/��/R�dd�pU)q,�+�y�Iͱ�J�Q�����p<�~!�� ��PHړ���(�דvOx���%5b��#�;��� Qe��Mk��ՏB~�����=�GdQ����w�� ��M���Z�kǞ{g	�7�D��9���Ҟσô�	�"]���'G+QA%��͊mn�|sm*�Lx���˺�ů�����[|����Ow���p)ǣ�o�(�p�L&� ��g�����as�q�#�	�o�H�Ԡ���]��jV�����vY���ŋ ���!��-r�'�Dv���$�I�O�ha-��W��t��3v|�e�p�3��!r vaR���N���6��һe/-���k��~���VT�)��ʱ������
��.j�ly��K�E��) ���^���l���m�h�#ߟ�����ث�!�'P6�-?���5�4��FcI����ڦ׍s"pN� 	@�	h� x��1�
Ȍb6�$ǳ�{�^S���5�w�x�/�ѐŝK�2��4t�+�ZG*�VU�`>�$3C�~ �KK��ו�J#a��ِ��k��B8�R.��6�	C���)>^��[����Y��
g6�h�ݱW����e[Ԍ���u�1�������p������h�M������%�>���'/��<�ӈ�E��ԧi��<�޷g�ջ���,@E�/P7��� ��3_�}%cu,�aJ����1��^�D�+�(�����R�X|�����.-���~�B�8k`�k����7}�M�������	�n�"�k�K����TGR;���m�����ɂ����OH��A�y�qPײ_*�,9��J&��)���bV�F�(�Y-q�j$b�A��dͅ��������K�W���� ��#�����"�<�'��Wt�0�N"ͨ%.  �V��c_����,^��bE_��Rq/� ��pڋ9)��"m��*���LR���H��V��`�#;1���W�l��$���$aR��1�6L<"/�c��*I��O6z�L�)��X��w,错'��.y��ř��v��	�����\^�##yF�X�X"��Z8��x
G� K��k�<\�u6���Wlе��,�D����k/:��kUs��W�ם�s�*� s�Jr���
�����0�O�`�p�q����Wa<��!��Vݓ�!i��NkĂ��Z<	�w��
���6��m]�1T2��������58�����ha��3�r�8�=��|h�x��aʍ	�F�ȧ��R:�H�������\�� ԕY;&��
qX��"��n�`�5SU�!P����L~n���5�������v4x_�<%BS�xD�,����孞,8����Wܟ���u�3�"������;�w�z��4X:�8i�xR�5R	4����'h
RŷD�ަe�V
4YWzH`9���:�T�*	lW��Z��]U�xN��mk���{č7�c�pI�����6h���� \Z��=�� ��/9g_~���|��V��71r��y�k>
]T׽ءe��m_\��۹3�*�e�[�y�5�u�>+��a����?��Ϋ'�Ձc��☕`����\,D1 �1h�����Vjm�����[j�<o�뗓t�jkxkSt?(<\�.�}�#.��c ��f<r�Iӳ�Io9��7L�J���Ǡv�����/sD�[�M�yC��2wt�"iY�#��j��I��Hp�|�C^�P�{
���X�� S���sQ3��g���yL2\��bwP�hu��F���Mh� `����P_\�o�����P�@9O�6���?T<���w����:md����P�G�?���.��u���@�G_�^�hR7|�����#����}_FX:�Xm��� �䞰g����2CxnY_��d9o���l
T,�(��ɂ�J[���y�c�SXY�0�g�u(uӋ�.�uR �g��у����H�k��t��ۏ� 2���x�t*+Q�G�[�Q��f��S�ϖ��S*�I��t�@���6�W��1"Ё�4A9�n
�iF�9
Nt��<��2rхH;�jo���)o���Q��+Ih�8_�ʮh����)������U��lo�`�1�:��V8�ٮ*�)���Ǎo�z 	��$Ȗ��Vd���
�Ѷ��6�~�}�2D	��P����\� ��I�@$��`��+�Y����H���n�Dv	�2�6�����{�\����'S0E�?W��B�=��24����U�Rw\�|K�����,Q��2��E�8����4s8�޽`�G�!smۉ�xu�2����g����b�M�͌kP#&3���ag�D�.X��-w[s[�!��P*��)�])��W�u�i�]?Uc�㹦u2Z�9ֳ�e�$��!҄]t��'�!,��\Z�a�
D	���>`��k[L˸��j�r?��F�Q4XN����vw�d�q4mT���۵�_�(u�������ZG1)g�E�^��
b$�sm��{W<�24e�.d%J�t�}o<eLO?�.�l��.���"�^ܖ�u����aKz F=)���D�{��������.�f<�ʡB_uy��������,��]A:o���N.�x͛?���YJ���DI2iAl y�W�����u�ә���C�� Ӟ.��	�Q�ö����5Y^�.��k<�5Puȟ���[�\�W�W�!�TB���(D�@��A�g��m���Y���n�vA��c�!β�n=Q7q^U�|n���A�E�|5*,��?�/~X� <m����j:�;>K��q����8��D3~&�"�&�J&�����j�3;��1�Ǉ�P$4�#�ԮY���rX�k/%��	 �j}����Ir�l� +����y�#����[b�5}�Z�1޷Xo��d2^����W�5$?fK��H֝M�jFB��s�1g�u#ܬ0�!Z�����y��&�C�p��?aOD���!g�=��!9�YDZKQ�c�H���*�h{n�4�,������X��9���zK�U-����U�e�������r6�S}?,�=}��Լ����0�XХ(��[�
m�Gwdg������[9AJ��Q�%.W�Mi�|����'E�B�B���f�LD��&��J�Z;�H˛Vڷ�I��~�8v�t���(���d�ʴ�s��O$��N�z�Q،⹁�W����L�׼�E�_���%��2~�
����� La�b,ݕ�N?t�6͟�6��ڰ6W�[-#󒕘&]��-��3e�,(OG�L7��z�eǴ�������AZ�>Q��+kضR�=�R�o�M��&���:O]R�Z?��(W�e�$iJ���/"�_��I�qxt���+U�[���c?�7x0�󢽥�A�jQ&�Y�b{M�/Z��cݗӱ�s��Ǐ�+,Q��[?&!��p�hJ�vɌՑ��fh'��@d��2L3T��	}�`���@w�'������p��s�R��m�Fs8��b�+���ݝ��	���0#��`�i��v�&<~�o�A��M~�ʌ}�����6ێ�s̈!t��$���'����5ϏE)*>��CM���By� ���zц���~ቲ-v �H�|�ǬG�P�r�?�_G<��s���HW:V����+y��0(G��P(v�=�!���x��L\.� �I�m������Y��-G��TR94�'l�[=��:Q������3R�ۨĜi����e#��X&���=�E��>�5��S�����Tv�:*�#�
�Qc�v�䝑��SN�9��7�6!m��R��rζ������D6]�-I��h��
�Mu���2%}%���S��l�qa������`����5��6<VI����t��#s��='\���`�S��:9N �go3��؄Sn�����&��SEE��!���&_�Q4c����Ή-���Y�ף�QǞ?X�F�
T��A�a�N7Ȕ��nU2�Ÿ����|����w�D��� U��P���2 \qb6d�!���4g�	�~�n�v��'�5���X#�Y��p��D��r ��L����u��ڊ���@�����b����P=fB�zS1ɯ�Q��*��IH\EG*3/%�r�$�4*��ȵ�J��M�3X=�M��)�\v�0�5�����g�{��$�@��+=w�G;��Z!��=��c���8u-zI	}���>�ݫ*���S ���2����]�ÐD�z���S�|p�Jl�c��L��?�FYğU��H�92���jol}�����7Q�:x�T�^J�4���l������x!�G�O�i�&;�XU�����߿�ᓍ{��
��=dfդ*Ђ�Ç�L��(mz��U��x�uH3�arއ��}��/F�;�⭞H�K��
(�.��!�Ї�3��A�<�q�&����=!���9I%M
0��RQi"��Æn�
�s�?I��E��� ^�V��{1%�'V���d3{K����F�ڰz[d")Ԡ].��ΙV.}��~oWm�b��1�Q�s��[\y#��y�#�u@���SݚO
���|7�t��i8{�㏪�bQ"S�h��V�ef�G����P=�[U>�I��х�e��S_Z�/pJ�}ה�Ʃ�ǉ�o��	j?��t �t$:!���3t}��5_ӹ�)�$د7�v,Y���q7��I�,M��E�u���.W݈�C��[��"�aS�֡���/�=:�,�>��	���꼲:[,93����b�
�۔�	p6���_xN���ǘkG4�K*�ݯ�S���u���F;c��8y\M��;dƄ��橺��+��� έ�Ҕ��C�(V�F_�~:� ���j�d�����P���Y�_�*�3�p�x�O���#�r}�%��������L�� ����G�����d�~Y����"� ĥ��6�P���l<@
�%fػ�l���р�>9�Y8�*6-��@��6}�H����Jr;��Z_��܏#0�����/TvJ������-�A�Bs(���L��=4*�OPF�0+��&�d�L>����iܡ����պ�������{&!�cb�O�Or�9��Ҝ�.( �����i/�X��@��/�_'�*�$�B��I~��N"0,so�|��srw����_d$py˞��/EJ��AζZ	�}����Rj���*�&��DL;�N�Շ���^��u
�# O�y!���cĠŽl�+��+T
4�ᨵNY��3���L�QF宅C��~��W��,���~e;<s^�@�ꍯ(Ca���T.�Luw�c��1~�����'���#�YmDa�w�c����X��Ṟ�#���i(��vk�fODl8(TvR��	��H[$��oʵ�����N:�/�W�+�x����O����qX��۪t@��,�'71��i�}d���\y��,>�֐}�1�rf#�?�_s4��p��<�<��f�.f2��J�Z�&Hq�xU�9&�MQ ��yq%����Ǘ	�-����[��F�ګ�%4<�X)z�6�ˋ�L��T��4�ɀ{ɷ8߄0N9JMy?b�����w��z^2�jc���x
E�ꆳ��2jbg��{�U:N��I�M\U�3ңIv�ZzS���c>[M��ө�C,���I����W���<B�yl���㖱ߘ��B�� ����n��yu��yP#�Є���vvz�����W9P,7��`UK��E�IrNb������Uq�G�n�\݊=VC�IJ`��C��=��2v��NR�Dj!+�s�j�8_ _��Vj��%CeP	�1j�G%�;�N�D����4-��)��P#�K�7�.� ��X;����s���4ؐ�%��$*X��ilvN �k���ny�����Y?uU����ß��e��ڜ���(I.���{�U�T�'�����R�{t��5�m��e��5��=NF�%pB�נ���D&�ܭ�F(,�_���z-�^�	Q[�o�j���U��_�{��bD��fS�{�[_��:�vni>�'n��M m���M��@fj-;s�i� Q��O��3�Z������"�M������Mk�<4�c�v�����)$	z>Q�ubw��U�g�9i�6D)	�.ǀ�щ{�g�X3Ȓ���K�bU���(�JPm�(�,�>d��FȠ�PU@6�#mw[��zQ|���՞�
+W���}�ӡ56�Z��0�y��%�����۠vD�;6�JW��q��A�q_��Bw�	,�1��� ð�l2۔e�;]ͨ~AgƓ^�!����j\��j�#}�0tXW�$�j����O~2��iV�_���|����{#��L����f�\� )^ZN�0�g���a�j�o�]�N�<��䆸����1�M=Lx�obZ�8]��z�t����X�1�N�P��ڞ%囥�S���Cյ`
�V-4(�O�ô�Q���쑇8����{�Vx{~��/�?_ױ��&�n#5���<�*�AT^R
�+���W/���ۂ�~C���/*�"P���K��3��+�1/�w�����*�||756�{]�Z��ܢӡ۽�#��D�(w9���ur��<@��y�����%�z=+�ne��1i2$a�>BaԍM�h������+��y������|�$������/� *S�VEj�|bq�R�[�f)R���䝩i)�ū�-�O�ou]q,3�t1D����'��MU�����2Ő5/R@{p��B����%�I��tg2����i�d���aW�B����p�RS�Pa�� U+�ݺH&�@ʏ�"0
��������\^���pH&ĭ����G�S1*�P�*�������P�9i�8��؁�a�9"O&��e�R��B�X)�>�����'y����Η� +$�`!��<�8�J1=ָg޳��u|/7[�����T`z6[�J+��=��s
�ִTe~��hy5af�����z��]���{pL蛌R��,���Y�Q���~��p�*V����dٷr.mm��Z.i�DX;�I��T��wǍq%��S:��@��]|8�\-ͨ�E��N�Rz���~완���s_	@��� ������Ha���j�l�N��G>[?�)���	��WR����������Q�J4�_��&-���ו�dG��̖К���D:(�t8JP( �<��c&nn�ޭ�g���^N��-���Lv�"��m���W-���ti2���d~��_. �GR����X�l�;� Y��za�D�I�ʺ�VW'"�m��k^��]'�U�E����ݰ��^��@)���+>g�^�%�Q�������#����?Sퟫ����z���EGyh �>�tH[i����B�odF���Kl�(!����E��)�CEU�{_Zٟi���ZA��2fbͱl����e?��S�g����uCG���ү� |4jO�#�:XoԳ���B��"��D(�������=���NR�Q��. h�I"��%x��s�:d�*b��%9]%x9��$��*+{�ñ�����hF �_Dc�Ұ�x�h@,��<!�����)�M�粎�г3��pt��6e�����F�;��2"��FU�̨���-���wA������0z��=��,|>���k�-��n3
�5��@W�j;��] �<ϵٰ��m�w^�)_ބL��+���	���Y�:j�b�F� �:?��5O�-�2C���yP��5�ߴ(��Slrl?�K����\ ��-�V	PC�L���M����O����q�b�D=f��.C�/�KSn�@T����-��g��D&��Ƥa:S�9�
v\>�x�T�#�L&`���SLa�H��L���\Q�B������&7nV~6nG���=ц�{���4r�3���s�#���=�ݍNq��,
\�g敩���N=F���׉=���8�8�����DA,{�E�A��~�C"w���N^��b�k�o��~�ʛ {P���6Dn�_��H���Ҽ\�=1���؝|�:�F��)�Y����?/5A) ������⴦̨[�'������%8v+��S�}�>�G*}el�Y*6f�����Ov�v��ʉ��;��2�e�7�{�W�_3/��QCgB�m�g2I\)�'��M��ir
0\MS��砆OD.�G����J�b�.$��^%�w�|Q�.�a�m�[_�>%&1#ǘ��k��863`6�\\&�N�E>.~	��5�%C8㘖���4g�J�׏��Ѡ.8���a+S� A���Ҭm8œ�/�'�L�#�k�O�P�(�+ʐ?^9o;arU��d�a~t�ݜ��{��Q"گ1�32�����Uu| ��F68�UIі�&(Rލ�5~�1��N;�-��F���4V�n|P�T� ^zB�!�;T�iY�ݢa��ݥ�����	�և&�:n!e#X��+Ct�[�R����ϙ+�J3�:�SU�} ك�EǶ�ҳ���PxUR$�����3�;����f�Ui�� ���x�J��z
|K/�O0���c��yhB/{�Y:l]I������K����0��-�v�̌=f�_2ӸZby���!�V�x.��+NW�"���
/>[��M!enb
�|�l�z�n��]�v���׭J�ƞ��l�Ns}J�#���w�15'�#�o�X�����Yng$�	�m�*]q�]�=�!맢��NF��:�	
���\bj���`�~��+w�R��b[d�Z�D)W=v�����XM���B�(]�sl`�m����Sq/�]%x*��lusr���@�),k��E\%���&m�������׽��TZCtY�>=�O��iD�˟|"���g�'=��[F�vT�w5�M�K������|
��&?�����^�J����"X'm�κܛ�jI�eA��s�ݘ�CTO'����%4�y��l8/McVU=?�G�كBp��e��Tgb�tY��el_X  /�`8��
ĺ<�
��T�
�� ��?�@4m�;�M\W�׋�A=�*,��x��x�āW����r�/��>V�DjM,7KX��)�d�d�
�s`�+y>ĸ�@q<,����16S���S��?nj*�����s�*��e������|h@�o�#i�	\N�k2���eQ|%L-x�J�^2~��:��:������Zr�V��ۅ�of�����VT�)x|�9f�c�ɰ(dR������\3�΢ͧӸ�/�x�5JHdޚ�w��0{�ﭜ�|��x�HO���L"23āŉA1i�RB@c逺��{mgh����4�`�L@�wR]�վ����|9������$�t����)��h4�U2v����K.��t������p�����aXf�a�Ѳc���b.�K$��^{�t�p}{6�����z�'��= m�r��%U��b�X�8c�f}1r����_[����@��T��+�_��������������D��AS�X��2 �m�O:�h��~�5��\X���a��MO/�>JҺ�(g�ɠ̥P����"�c`d_	���U<_�j?]HZ���ɺ��8x
��d��F��ϫ��j��_|�'W�����-;�T�b��Ypn��:��*1(q����c��&����Xr� |���^ �i���G}jB���8@�BP
?��J�P �`�~R�$xm�x���D�����W�s���PH�����������߿)*-�u#t�/��su�:/_?�����������>:ն���)���Ĩ�O6�q}N3
9������8��m`hV��1�&	+
j�Ż�;.4/�+�����W�
EF��O*�%Ď��n�Zc�K�MX��貂�/�9�Ad�U��"�OCMn�_-���5	^K�3\���#Kإ���ֽ�lk����wZx�K�2�h	�s9YmNOC�N��5S8S��y���DTY�hR��NY�k�����oi�{u���Q�\u���)9���X�%"05����9:g`N�V���>���T��J7��AS5�	 _��"��6�p�����0۱���սT4{��UD�����ׁ�5�D���F/���,B�	��HOb��d�w�!K�"*��Vx�}4��R�׆#̈́��W��.�B��
���Eί��u!��\��
%��(���@�}J�ŷB� �;�"S�������	���n��K�L� p¹�ҠX=�T9�>�F��P�0VV�Xj�X����.#�Ͳ���mQ>�IT�k�����(w�8Q��H��2Xy�����/���e]���
�w�Λ��a�ͻZ:��ᕸ@���¾��"��������;s㍋0�z'$����7^Ɇf�((���)&w�ؑKJt�7L�J1V��"�x0и��������; ��f}x�i=u��t���?Q�$(NJp�G)�t*bȌw܏M�jXN��L���Qϐ_PU�;o7��x�(��*�O�ռALR�B�3��.�r�σ���]w2����c��	�(�w�����dӡ)E�O.�V�M���=u�i��r�L��l A��Z��+`������١F��b��WX,ŷ����{uG������a�"��$�V��u���g��ޓx�k�Y��+��3��"��B��h�&��ҩ�tǂ��m�4V� s�M�i��W�I����e	+ve��[�.��lyٔ��A����PQ.����*��"���4種��ު�����a�$�NB<{0B�"�K����ES���W��*3��
��|ڷ�Tc��
�C��K�-�?Y�����3E<O�����7���/�w)�;�m�c�b��ۇ��^op��y�`;�~�H�,*�M�s�i�L��P�Լ$+@8n�I~<l��cu��8���J"h�+�u�B�$\B�7ć4���P�('t�g窏�ur��%ʲ(�+a�/Z����S
�w(x�Bv�io�a�� ���^l���oGd�Io�(���B���v`X���K�ϧ.fHH���L�b ��e�
GW�h�8�D���yr��1
�� U�X��D�R���l�W�[��'^��<�(��B���R�D2@:Lt�Q�(��;�c��t^*,͢3�E���; e$��Ċ��'y~���#���=t��lغ&���}_����x;�sq����²�l���%����[��S['�0p�pٟT:9֘�U�i'����ۧ�ߒd�
Qdە�i�S���n������@z���Y���6���>��b`�����
��?�}k��� ���
uv�A��K������望�}of����	�Uڠ|I���y����Z#�_v���'zX�V%s>��|��^�
������@�X8ߡ9�SR��������c�V>[]�Dna��r�S)5D_�۽�k���;�N.�>
Y�x䲋�-�K�x������0� |o�jkd0eJ)#�.��T�Jq�&sI+a�m h�iZ��fo5����1{b�H?ߊP�wU�7�K�������N�!Q���\��~w�e�N��MN�59�aʯ�\�T$!z��Z�����*�v�I2/W�o/��'*��t\H���8�ru�� ˖ Rs-B9ȡ��r��AK����5�݁�1U�|dw�F�."��*���acS�Gt���
�ߧ������2�u��yj��_�������x�a �p�S���@q f�������#��9��b�+��Dkg����-��sǙy�L���c ����̨��HHc���7bi'�,���L��K�J2e�b�֧{lfo�Kx캙ټպ��ˎ��.Τi:���A�֐��eeoXW�+�	�06��|�bl�T��[q�&S+��d�@���Fd�]f)5�X�?�j':}�-���G��Se���EH���*N�R��Q���=i�$��A~
V�-�\@#DHd��D�rU�Y���~1ot2���x�oLǺ@�ϭ� ���"�U}���P�k���ݍ���/��o<���S���?#�C�)G�BE�&.T;��^^�ų[��}��0l�7r�.�]Aj�ί�����J������)��N^�A��m^T8�q�J8{�P�G�Tnd<X�혿��N>gM%$���`�~�]�Z��*=KZ�!���m6��W�A>a�5�R:c6����d~*S�*�{[Z�|av煯��\��T�W���~�J5fK��GiaR+�c�e��}9�)'����ey�Ä���'�f~u�� ���U�@����C$��+8A�n��9!��	t?BN7���EP�an�f._$:�d�����x47��/M�͖��U5�C��v�{�h�)��$� Ϝr.��ѮO%�����,�����Ve���4O���b
R_Q��(i�߫��?~��&@��� �6�\M��QS�OmُaɛCtWQ��y���6ʝ&����*6�GO@F�����V�R��4N곗!�>%`�\p :N��\���T ��*�ϔ�D&L��9�A(�$:�I+n���M���=�q���ŝ��% �c�7�$j�Y�l����n<�$M�d�>��T�e[��%_��һ�9������� �R�!?�3	D��� �um�6`O�+���og�'�\z��A�[�O��{T�:�C���;�=���l�-;�9B��b������/>/^YSgF��3M�/� aY�!�geX����x��.{�y#��c�_��"y��^�6Q�ص:��aW��۷���ʣN*\�Ks��Wݳ��9�{�3�E\XČ�1�ţ���z���q�n�?ú*�&�Ɛ��x�Z6>�WX� ��M��o���%�C�f��@�}��(�P@���4e��sQ�W�iC\���f�Ey���1#Tj[[x�?{h[ݭAY��m���)A��(��Ѣ��r�Rf�xB.���V|�l{��%�G�d�@dł�&ϓ�0�0}q,^�F'���j֟�۫}i4��5�x�΁@G{E�7"�6�c�R8�~�����@\[���!��+�Lj��Ͳs���i�p���ML�c����k�(�j�����Za�Z�)@A��Ew˞�!r|]])UXL�;#NvD=3�E�F�By�%3q��' �;{I߷[Q�������/���h�8����.o�(T�59�����2p��B^�9�����(�Ѿ��4lK��\�uw�h=��JP�,N��P�yz$C[����F������y|�ɻt�g%�z{$*�S�gi�(ї	�+�n-h�<UQK*�tǯ?@�u��N��
��U��&	NB���g��]N֝�n"���_OkW]j��>��̠��b���}twa���O��0���1a,1e ܶ۝�pf0Vw�JuR�^�WF� |�&�6|�Z�f�^>�9�mb��j_&5F�v]]�6�2��,`���h9�I�uyG��E��יqA��G<�Ɵ�}h[P�~/ל'&6�g��J��Jm���'LnLD�����c�E�3�H"�}�ԺpZ��UF6�<-����04�/U��!���>D� b �%b���o��k��Գa�7�����t
�պ�l�Ș���!۬��g�A��X����J$�
_^�T�֓�6&�QK�\YוSQ�z�Z��3�WH����l|�X1u�Z�H|�L��H�ʗ_k�� W[�C¢Gi7�� �rG:�$��!��W��3}�G�{r�w�W�< ���c-5�Xq;a15xm�0��+�� �-F�� @�	S�Øo*�l6w���%N���C��-��r������hÀ�`f�.��,In�b�A��9��k�2���J��Q��9J���0k�B���Õ�#��\D�r^xl2&"�����şA�)�k,�Y�و����&f��x=��� ij!���;y���o�Nm[��0Ѱ_��-��Ey��f}:%���X~@p�b�GS��4�	SHWd��]>�:R��.�P���iLη��T����L-��_a�l�9�(���ɏ�$�k��W�����?|�-WM���p�S��A_�}���QQ��:���:fs\��ބ���u����䢢g��ھ݅2�+�Z�3��W�2�q�B�:o�2ns:�dM�ړ��Y;L��m�PF�(P��'dߠt�PMyZ}��h�"�eR@.V���5� �=��"Ϭ:-�:����^^�z��Wއ�d����Qy?�\�)b�	ϭ^�^�q�fI-���~��;*���Zɼ��g�3|�n���\!��i�U�X)��@����t�!�)�^�� �g�7j`��\�9�zO�s'�?r���q�I[F?6��R\�*��;���������+��Btꎹ=�X�	疥4���v��Q7?�j�^<H�]��Thv�&� i&����ڍҋ��^/ǝ�F���!e5��K��2��#7ލʨ�H(�א �2�>��j�+D>��STܵ����A(
��yX�YҤ�%~�����)>��ũ��2	W�	.öCo�٘����	/�D�����!-�)6]����2�!-�*�r �V�y��6,��.�P��3X�S��0:ĶS��)�o���E:�D�blk�SY+^��$���ۤ�����X�/�02Y�ǡ[�ZDnW��cg�F1���X��-^%�N��i���A;H�q�gؓ[�=k��j �~��Do� <M����:r�<�����]�%%Ye��"�i`�"���Q��&t�o9v_g��)}�����ҭ#=%/��z�%"ťg������.�L�)�S3�C�1c����Q!l�=��~蔞ܤ����ەq?�8+���'��4�i��h�a0^� q{p�i���p�s�;J�S�v{�ӈ��c�W,�d�D�+K��4?4�\�G��ck0"�r�����hV*�Xzg�s�5�y+��i�Q:tyP�)�����ŷड़���\�D�. o�� >��0��G�����05mψ�4v���H���'z�ݾ�RD�Շ�\ue�Ba�vN�;�(�C��׊�z�՗A�����O٢��( 7���\5��k^᭨5��=͓CK?��p���EQ_���`�&@�4&X��2�9<RQ���$~���2�9��$M�9
�Jf�E.W�P���8^��lЈ�6��4����S���,,��i�ܚ�R��梓�kg�����ٗ2�>��z�	���|e(���4��ic�Y ��Ym����1�X&#&9-��5 X�
��6�@al<�,�I��]�����~=3��Z �����w���;��^0������	{�2�Yꥩ��7|��2�S�e�����z�F��|y
��\��w�)��M^�̬��h9#*�~����xֺ�M�Fp%��TPfפ�tL���>�=��$�Mx�B����U��6t���{��U��`d�{��f/�31���s���j0jVߔ�L,Z��2���~������M�*�l���fG�2��u;�B"k�>��q �~S i�P��u���CU�hXx�r�y �U(4�d� Rr	Ӄ|�ERQY\B�j�i�"�P��H�ْn
�3�]�ڀ��YԤ;|WYc�6k9-�kA��D��*�8�&�%^~v+=.9��#�GP�"�`Y�N�C�m����5Ḑ��u@�B[Ve�˨]e���ޣ�B�ʍkԉP��k�^�Q��P���#����sL+�/�}�A�f��8~Q��c�=����+�wD�*��M���n.4TL��t��x�����r�c�o�}I敒��4��0�T��9���T<��*���;�я*����7=$E�f�H���l\������&���Lp�|��)a����P��]�������D�brA�ՙ��N���^�ō\=h�UI��� �<t����������_�H7��ql���PO��M%tXӭF��9ߒ*�1	3\pnA	�2��q�8�.�OY��c;V6������h��Q������$G��T�}e1���lv�S\�����{�4����J>�/����#Ù�Q���ID�8�s8�彝���O�-�+%"��6r[.-��5��T��R�F̦�RY�}�K�ڑ�8e������ �Qܐ���U#@�%�V9�O_>"����Mo��p#��N���Mǣ��}	&a��Ib�,���B�3SA
k+�?��$K��zݘ]d	��y+�k�"��:ie�j<�v��TRP�0��c����6�y�����sG�ajC��I�>��D{,�% ]�0WC�o��0p�{QG�~T��U�6df�Mv��x���z���e�`�8z46�z�E��_���s��h�6q�:y��aA?��n:��Tmq�%D��z~Rw:3#u2�n#��膹u9��P���n� 9>SZ2X�EMTewm������U=�0�$�8�p@�O��4�W������:Fl%_��3'h��7�l=���;C�m5U�e�����G8��H/��3h���&#���&Uu�8u��[S8Mr�.����.aD�!��a���?�m����>+�]@�?�$�o���`�x������'�n&j�͕#������@VC1�k�9�e�9 ��D��P���B6�5xЧ)f�^�[�<3>F���g�L�Ǐˀc/�O�M.��C�Dq׼$��&���S"*���a��qD[p}��7�/���֧o���r��"{���2qGr�<2��2�ۛS�X�pC�.�։�8��7��"�#��#Mpe=h�{��o���n�G0�0H�Z���C��u$e2t��F��C�[L�sT�7�?���?���s"bޥe*��{o�[-9ٻ�5��~�>�c�
�;U(�/F��2�R"��4��	qg�fU�Jޫ`�:�Zb}75D��qE����#���Sc>e<�^�`����@:}�UUiۣG���~�"0�����)��ڎ�vL9��"��9�Pר���^f�d!���$�Ҫ�D$�j�s������eϟmB���|�^
�Ul��[
�{��@��4v���|�N�D�?~�AQ������~����S��±�����]#���vrGh�-�Fx���	���X!̟�&�Ú��a�~GJ<aʨ/�ɍ)4?����x"H�����|n�O�#����8d��`�����=.Ѵ����'D���#����H��n%��e�#�1-�M�CA��&r�Y�+�������)Ǫ� r�T��*{{5:%D������YZK�>��)Yh	�nu����!���/��)  (�^��2�_v=5l|T�Yі�Wn"�t����W.�n���
MYj7�|^��-��]�Ż�U���`�L��u�n>�cJ��y�#��S�2~��X�r?��Ҧ6�!e��O�x�&1J�����V����m97�L���zy��"�b�Lģ�B��R��X��H��G>[V��n+��oqex���4l�1T��| ���UG�i���,�C\����*A�2~v8pt�{g�]�E�7䃻��(�ɇ�U��5Fz�@W�d�݋K���t1U�f�$�m֑���5a�פ�����_n��=y��0M�Q�r�����{/D��ʷVK�6d�#"s�+�R&R���3��w�º�	z�1��\���BΏ��d�c�/k�e��	V�"��h���߆�+��j�C��d��g�jC�|���B>8X��ހ���G� �'.��c�piiK���26 �Lֳu%�#Z���3A4��.�u����3k�T�~�G�;�6Dq ����UW�J�z{������Q~��3gD��1E4��e��4%`����R	�}o7���g�h 1�����3a����H�vR�)��.Ij�^��M�8��$i�:>���D2�~o��X �R�\2��Cg���WɃ�%u3	�>}i��y���'T~��6�(r��;����׬G&��6�����wW�����2
.-��,��'v�#��wZ��ZeBپŢ��Ƭ��f,4���gx�i�H!��uΉ�+q����g��?�J�3�*��l��7��e����a�I0uٗ�W,�CV���;X�Vn�qJi�.��w���|�Ǌ�~���	6��zb-�&��[.��sTw('���l�n�h���9\�0A�=SB���<3�N�<�?|O���?��	/��U�e� �����P�=%b�����|�%�D��P�e� ��<
��1y��{!��+�Y=�'e��5�p�l�i[�/,�U_��n�Tv����� �k���m��3�϶�)03K�tP֯�,�Y�>N�j�s�xLڞ�#���Ɋ,��Nv��	h;� 7�#��m%�ҪJ�C@mM�=z;�^e�_�}ժ}0
�Zx�VAZ��ơ5��U��u^:���wo�����OV�(>������M��u"���,�wnd�/IA4��1>��b����NX�YH��"����ۗx�vB�󾲠;�z��Z=�&��	��1��(O�5�4;{�E�T�v|X��}�ktxO�N�+���ԩnw*��زc?� 9uۤ�&\P�R���&��G�������?��kuϳGX-j�"b�]��`kO�uxù�z���7�XÚ��v�6�q��=>�6��͓��i���Ϧ�*��x����z�p���:х_�t�,pj�t�j�+��t8U�2��b��"��\֗�f;QI8��f�qԑ?��RcM���O�����ܹ7>�w)�*C�,m��iK�/ML�5����O%ܓy�4fI0���~R��2P�Y�PA39V ��/Y�%��!�q�I4��{Gh'��%L�XE-������t.�,
��wt����G��/p�<�1%Iz���@��ҡ��l�����c@�h����0L�V_&�8c:)u"���+�6����w[��R��l
edo�i�B
�g��!�O��x'��8�9WWkٹn�O܁��;�����xF��+�Gn���n*3�Ѳa7,��)s�`8f��p�y�b���
B� ������9Ȝ�@T����r�^��P{�����Bd21I��s� �b�{�$��Q�t�x���?a$�
J�jf�]�߭��>)5Vi�Qڸ�ml0�K(:/������c{�1���3�����S>��Q�l�!���ȟ�Y��ɷN�2���f�<G�O�jè���9�&mI�{qJ?���.ۯ��+h/��D�O��%�&�51(��ު>��e�W�D�� H�P�8��82��%`�r�����-]�A��l8�KF�d������Ya"���t��g�t�˵v1�3�w?7/�>�3�~N�O�3�)���D]�2���O��j��,D�=�к6s�P��>�X�����/���܄�p �&ҫ)ت���	������{ɥ��}���}�Mue��f�8i�[ �7g+�=���K�ݛ��}� �Y�u)]8qb��ڟ�Z�����U־��YL�vj �6z���!��h�X��@/C����ΝΒ������� ��AR�r��o\ �O�`��M/��ݲ%�_S���>���ް�(�?��*�����(׏C�y�{�Y��B4O��e��˪��by�	����Hp}��3U����c�p�J�5�7vl���%w?Kٷ�uqkp��Zh��/�^MU�.ؽ����D��(8�Vy����r:�ğ߯�������!
|+��I��-W��Ƚ�5qV���չ�@E���!C���-�c��N�ߍ��ρL�|(�ʃ��VՏb+)#Q�Ⱦ�v��i��B�et�{j���k��c?�$C�]51�N�]PHU�`�r�5%@��ՈP�MT��&�;���!,�֯K�aZ�\1�>x��}���P](��,�Ц��t���<y�>��������[]�s�=
�/a">g�`�M@*+^��5���mP �[�U�ξv�IzC�f�X�%E։��ӫݺtͮ9�:x��ܯl#�0!|Ls�a}/��>T;�"?�c�x~d�p���j�iV8�d��0t?��A	@j\wI5N���@���\��� ���[ ޻lN�58i��hY^�c��u�6�d��~�_yY�BD�˲F����;y��)�(EtĨ�~<T>��2/��B{?���F}�$�Q������� -��X�F��������F�L"�I~XYI��ʙ�<,���8�MA:�$4����6RN0P2y�=c��H�y�'�l�Ȯ,��aWH�F�#��Y�Sˠ�e��@	���~#�,<���A���M0�y��aQ���r�XR7�n�$�'���U�߯��|XKzb����̈~�U�,�bO>w�J���ќx,�e��}j*Q�����1�����_�҇a9�VJ�>�15"���O��a��_cF吥WZ#כMw5�R�5ar_�E�*5�r�嬶Ӿ��⡮)r��O�K�;�0H�X��p��v��;���[q�;�9"OvA� Tg@�nO�=�8Ù�$G���(����i�Tc������?�IZu�9~�\	�h�˨d��)���*����P��y<��iɡ��]M���gK^.�;:��V�D"�?��}�9H9�6i<�t�����TJ�N��F0�y�i������fE7�浨p}\k5G���Z_*�%�Z�9yW�@4ِ:ߜٱ���v��z�q@2/B*��2iD� �Z��Z1����	[T�r\C�d!�SѢ��t_X_&	�<z�fc&P��;jI��u͔ ��	T
#~�����f��4Y�(����:�������I���Y�Ǯ��y�_��S`�
��I��=�f~ǅ!���#���} ]���7����[����
�XC%�m9A �C��Z2.�Q���x��K�P*�.�uqG7��6����SG�Κ:��6���%$�s����7���ʇ/ȫ�+�`�V�j9Q �<cc[Q`X6�&�,����y{S����s��Z��dWU��V�)$L��5�B%&����4�������"%�.WJ�	�E���09�=SA�8Ca�nx4�/B��nv�]�֎h��>����^y�7�����Ϻ \���*������qev�y��<�&QS��|HZ��Re=��?���"I�F�~�8b�@�J��n]8v��`��aҐ�o
2)��ֽ���Q �l��K	���:/���������IԈkR¥�� "���xݰ�gs�f�I��j��=����(��|�;�MAdu�t�m����ɳ�sޜ��2s�Y�6�+�"���Ժ�;�b�Q�ϢB�wo�;&�ȍ� W�K-g���K�қ��M�0�먼`5��� ��9a�Z�K)����E�=S�Y�c"�P�;Xy���罜>��&�	3M5�I�of:=�J�m��֌k]�����J?>���K�e��(G�C�H�Bj>���`����I�~h�MX��7�>��M2>�/�7����!)�L6���I�ӞXx $�;4�K�Ly��_P�5���t�OT�L~CJC�ƌ��ܠH�����&�>U�5������
�& WR����9� ���!%�n2��|�~ �T�7|�@�4`�`}�����Q���{�M�,qC����7��zN�.p�3ﶿ�N�+�� �r�v���Ej}�����G���R���:+�q��ING�	@�nwsL/��7r�jj���(k.�$�c������re�摴0��=mq>��Ĉ𯑑�8'w�̕�Ք��^y I��c&<�U��}�1�qDB$�؆t�}W����G������h����x�Qu�}����Ne�ӗ���a8�oW�d+X�Cf�w��ev�[jE@����i��Gt�o�)@X��\�g*ԍ�����Qf�⥹�&.��~s���g�Mu׃@|�/#�V.w����8�� �H���Zp��~c�s9o��5�yB��^��E��	j�B��ǚ�3��~�z-�����)��g�MQmp�/�j��0�qT�B��F��^��e|���9�l(�
⬛"����_CZߔ)�o��s���@��Odz,���Y_���g)rfiY @�� :����k2��0e�rX�4��*ad݁7+���u����]Һ�DI��3Ax���M���P�
`s_���E=�Ĳ�+Z���yG�O�ʂ.c^�u�Y���=���ӑ����ok�d�x��xwDQ���LV5D̥T�ȣJ�/��,�nڭ��i,��L�'�LL �n&�qL�� �Ȯ5��%��欙���[��ί�Y�W+��h��k*.8IiPB�[��fe�{��"�R�����Lp�^�BL�C������	�))��>�.>��� $�7����~C�e>��m�X�^�bF��vÃ��0Ԋ��|k>��[��A}I��GC�K+�	S��o]tC���������ԇ[G�g��G�A�e��vYH�1~~�_�4��hW]��T�Z� p�$>�aR�)ދc�%L�U��T�ک�����ÿ��Eޮ�=5�F��4�r��b����*�S��<cA6K��4���6۩�fᰈ�݆FN�*eG)rna��ǯk̈́���Ā!	�����|�����t2M-�3N���?�%���"m2�.�����Rb��@�S����Qn���Z�fM{�6A��`�>4�8�|�]�
���16���?0������\q��iC%:��RYw25D}&�f��h�=NwX�5��lÄ���K[�O������F���F\`��{�TmN:�� q��p
��n�?2B�H�Wøɕ��ͧ��Hy���XX�� \��L/��?��ع����|�E��*�5|�͎jh�f��>J����,�:����a����H�7@c<'�ȃ525r���'�݁m&���/h���uI���>xƴ�E���cޥ�$%������45Ԑ`0�j't���-�I�{4b�
,޺ׯ�C���F'�"��|[x�n�<_�(I3�P-oUoX��J�xa)u^ȕ_����'�{�V������_�+=�4�`�z�N�4ۥ��%Mnj�h��P������X��[Wea]���r�M�ī���q��qY؇�5	�q��5N�m�XF�j� x fA�2뢈9�-�_ţS�`�8fU��3D?y�[���{���	�M���-�zP�H����۪�I
���c���Tɢ���o����Ǽ���B+7��ӐiҖ܄���=0��/_>Z��h����Q� 12a诫e��^��?�;�v~mZ	��p�tC�{�I.�;�c���<0���G�!���{��ʞk�G!�n���������[Ʊ��pl�i;h����}�����8^PM17ݺ�VAZ�����YB�\�p؟��^��%��창U�o�z�����q�b��k�{��ӷ���6���[w=$�VC�8�?�ۜ2K���@��țJ �T�)����Z�bU�S4�S���U���c���������5-���� 2�Sr�r�jnk���~��܍�'ť��tc�24�T�ٸ���E߶a�}v�ȟ��e�T�5DK���ҕ�J�:Z��6�_�%e����L��/`�#D%�At7�k�U�+7��J�=�F_"��I���؋N�/k=
L�^���c	�n]�	�Q_��Ү`XcA�.��K��� �֩�k}u#Mv�M��51��p�"O�ɱc��$P`?4W�\��~E^ubn'R��9��	?ট�"��T_f[�m�~�m}�@I4䍙�z�^�ة���!�h����Ǚ�$�'Yz��AGlM!	)
�o��Dؓ$A��T�Ɂ7�C%^���qG���5�9��#�CQGC,�4�au�7��XVe����o�^?�[���~��lu�:��˱�#7�f����V���a$R�
n6ɿ:C����\ɺ�CXɎ2��+�i�K ����񥹝�~ʫ���`�t�[���%��P'D�4c�{��.��1"�hj,�nh��Wʺ��,��,B��:�4���j�t�I�.�P�'.�����	&_����1���Z����n�	�_&~6��--vk�k�Fx�t3`��E�E�xj��/|wt��S���YE>�k��R�F�,�a%j�,..0�m&E���r��!���e
b��GŔB������6_�RSZ��:���܈�+�Y��4�������oٺ��E��G�c���Ly~��郵�qJ�ث.����f��BYk�.�_wNkz���-������2+�$�4Ţ�g�y5o��r'�O��Gh7MA��*J�����'<�7��o��ً�n��Q�85{W��&��
�mXT�;zd��T�m Aq�eJ"������0�~` p�JI�����%�d�1����'o������B�m���>O���NJ.�KF�	���(�k���,��?!F����.�d�1y��`��0���\�L��C�+3 d ��j��yq����던D\����
"3�T���B��'|m��!X�M�8�����o����K��/N`�m��{Y�7�H�&ż�,z)�Wu`p���w+�z`{�Uuل#;�81�r�����{�Ar���Y�M�#ȡ�|�U���\����ϊ�4�#�~��ⴈ���P�v�m�򡸑����"ZS�7z��2rZ�`J� t���f�)�#�6��$]0�=׎f���1�c�-@���AI�ܵA]������y�K���}q�q���?��p�o\}�@~ݭq�%�Fj�'�C)��!��,��)���`@�&�{E�hs2��y?����vZ&����(� �9�Yv���Hu-�����m����B:j�;�CA�<|yo�H������*���#�%�Y# e2' [M������<�>�s�����ɰ�����ڴE�.�߃�{�V���U�[9��`��"A�v2l����/R����p�[h��K�
�Ԍ�DD�G�S��J�&.���&BC�f�ؖ|��P� ���/s��~���\�Tk]�Ւ
l����^���e��m4��;�n�2�D�9����R����>:���O�Oey�T����Fn	����Ć��"���]�	�_�qLn�yI��	�i=y��&1-�O��M��h¦����� s�+�?H����g3��A��@�{����5��:�Q�� ¡�,��n���մ�pL�۹J+�^�iy����<�T�/����6;��m0��]�L0��X+)(�%�l�I�Y)p	��n a�$U��g���v[��u�e?W�q�ȝ�]3vw`��Ɖ�t��Sr�=��J�4����'�x�歬_	�N�+��2 ݪ��_d��;���[L�ܘ5�Ed vY�T�D&M�d��r	O�C-C�pVQ����,�j���%c�cdb���1��U(��hY��r�'�Ps�5��h_�e�"|�~Rv��`{ ���ˈ�wm���:Hu!k%t��̩nO�LM�]�*��X��q��a_M�RJY<�a�|AT��gaD�z-&�bd"|� �~�{)� �1GfGՐ�zխ'J�Gד] V����$�[��ŦtA9cj��tQ�Pal�-��w�\	�#_^@���k*���(��+7*{L�����A0e4�3~J��|��z+'C��1�a����H�����B\$��ՌHF���x�x���o���~��hO��-։�$�g<�qJ�[�D��V�ͼυ�sB��~ᒯ�D�2���N�����z��g�Z��Q.�=�6�dt�dc�'�8�=�II�،�,�Hۋ��dS��:��2?�<�z�)�q��/�Ҹq�!h�QV���I��-�2�ǋC�sǌ���NOյ��hA�}���a�X�C2ַp=�)r�/F��A"I��3����[�M]���H����o���"p�n/�aa/�z����ę���| ʤ�/�_hò���F���%ޓDD�V��x��;$�J�U�CH�%\;��}a�ū�Gy&�BmF]�ي�&��>�O�8t��Ƥ4n
��*�Q��}�H��>e��`%/�IL��>��)�Cp�l�y9��ܨ���Ҭ`�
?�k[w2B`iz��گ���Ĉ{���8W�nW�G�NTgM7j#L��qʪ8r��*,�6/�j[��V�p?Z{~9%�u�Jw�fJ�Oʎ��R	����x�N��q��#Uu<��)����q�#���é� 7XW<¸���-�&n?���]E�p�R��!K��<��^��w#sYp�揷��h@rbC=nF*�����{�B=7��1p<���	�o�c�u������r�B�O'�K��N��`;Q����m?kh2d�����?���9J�B�����:�"UQ���ከ�j���T�0�2��Y��bq��~n� �����X3^G�T�B�(`q��B̪����������zOӊW��j��Ki��i�@Oy�����Sd�m{i�u/s_$��	��Ģ�yy0��Z�DQ�K=[ �X�b����j��c�Ԙ'�P#AѠn�q�c�����z:a��BK[�z䭛�mD��:�@'�2���A�y�,D
��k�I�p�����\������x��A���Z�z,��\Zo���=E��Lb)
9gԃ,�Z��=�zI{<hz��ÝBMof��!���j1&V�R+0*����ҕJ�G�R��M��'����Pv��c�"��-[7,�^&߲��_���#d&P�t�y�⺕�V�dZ�jc,���4�{Y%,��#��N���h����hƹ!;��j���튌'�0�����!z�����G�b*s�Sȑ�Kz�4�E'������q�j�D�7w�>�-�-١��E��R Ũo���̊��yh{�&e��4d��` ̚a�	;�L)%T$h;֫ڝ���Ѿ�MEX6
�m�.܄�KV �IAƕf�Z�w�b�s�x�����y�͟Y�S�������`�Cl��#���"��'[�,L	�w�J\3��U^6J�<��6���l._��/l���5��oA�4wFps����ND��!7�&a�Q������[VA�H��@��E���ҡ��VK�Yr|��E�?�/�����t@C��I�XU�h�����2߮���͈OWh���a����B.�T��!0,�`�~ϵ�b	�Y�Ș=J��
P��f��qŒn�������A���U%��"X����g�
�|vmc��Ř�~we���|3����� u��U DWx��LE��Z�������O9��6�9dp�h��y��������)md�G��p���$k��z�������������(��<��@��76X[z7�=/,~|����<��)P�J����r,:� +M�/,�\0�[[�� Uv7-��zP ��s�	�{�ĳ-�I��η��I��*�01�51��'��]����y*VZ�SuǏI���������&obP8.%���C�@�[�K㞏UZ�s?ڋa�U}��~�5��%{���%U�tI�lN�In�R����W�5 ��e��z��T��x���"t+�*Pk'�?9�So{�|ܗ$������������t�u?��#}}& ����/ ;�!6�	P{̐<p�6�0����Y�M��@!�V�ݗ���Z�+�a@�\@�j�d��h	}}uC3��K�#>�'�s�L�j �&��'��٤�'$A��3��GJ�ԝ�L')������ȐPt<?wW���h��� ��|/@H}�?���Y]v$�a�K ��o��]V�zӠδ�6��\���=��85��r'��I"�CH����"���qcMV?b�.����,D���~�d)�r_|kV3�-������%��"U��Rq���b�ј"d��8���{����3���[�E�5N /Y$��X�U��������4d�s˃oF� &���2���� 9��Zh�S?��o;���#"��'�XoOvH�Hͪƪ5�m�їq���/6�����w�@���fK�7Ӫt"��(3;T�!S���
q��Y�n�������Ai!��K&;=6B�_�:('e_4o�GL�-%��Li�ǝ�e�2;Vf�R���0�ΚS*�����Y� F�{ys��
h�aB[��(���Q�ݝ�͈M��.T8��x�.v'��g-���M�YY��}'t�� ���L�`�M�1,��{�$
�������r!Q��/������,�R��� t�?䟰�g�m�Ucn��r���|��c��/,|L4y��3�	 t𕗚7���`i�$	S���}P�7[�Mz��0�e-�R���@�1�J�g'qCٕ2G`n32ܤH��a=z y������ͪ�?�(���	�r����	*��~�h����G�0'/��R�kk \aN�Q�"�$63{o�oI �O�jN�?��Z��3�5��FTK�.̾���@D�5�20k7s5O�kj�zd���П ����e��rйKr��^�)�f��r���M��bg?��q�9f/�
���\��9���g�+�ߺs�M襨:��[����=v�A-b��^�
g�-��e�QQ����|�{�%����J���� �t��ϰ�'���8D�X��Љ�~VO Z���H�f�D�d~��vs��f��*���h�|4�	D��]=$�V4dİ���G�cU�S���;��i�lSN?zy	�j���G�4��jL�qs��Vy�W9���Y7�$!2	�ݯQ�0����qɥ�,��]���{�O{4�9�!B�����Ȝ�p���c��Hr#8kh���.��ϱ��5��?H�:I��)���6ؒ&���~�k2N�W*��]���s X.|��B�aB$�\r-�Z�a�͏g�7��t�%y�[�jB��a�T�2�JE}����6�Iζ�#����R8Lxae$ �8�cTS[@{�������H�pѽ�UO���Ƌ�����McWR�h��$C��"��]x�I�C�J��$l45 �bC�wN,�_Y��;��Pn�Y�ECSv^�1hҁ��IA&�r���?����r,Fa�i]��%BrZ�m"O%�PJ��?l۽�I�������<7*z5�Dc��Z���VGK�c���Q�<7�!�g:C�sW�7��hQb�׌�x�T�r������i8��1�ꯒ��٨�^k��$N{��,�\�!9۰ڙ�Y�i`�~X�<{pâͧ��ugwG�g�I�0�MטߔE��7=]��`rjG��F��0�� �%"'�nX���8w����Ei����]���r�,����/ɂ'����)(3`�0�NitP��.�t:��b�x�VOڂ��}�\�����	:��xS(������� f��޺V�+��{��m�y�x�q�A߉��NYwd
����A���#��4�)v▪�9��I�1��$��*p5&t�����;��ͺso�FR�Om�������C�_a��Qx��l�ˎ��{��0T;
Y!�K���7�XZ���9�N}:������ ��_=B�ע7�K���B9���#�;���V}�`��5yq�)�� �lG��l<4ht����v7zh-_���O�Q/�H�C*@:�
��1 մ=�K�7w��|/���RR��?����%��Z҆�d��b��'t+��Z�U�l��<�Ĕ�^!�a�P�p2N�J��(�(�f��>��Cֶ�aWd�W�[��`��y���7jK��ٶN|q�F���
�Q��X������%wv[��N.���F���� ��eG��}4h(�7��'ࠆ,����?J@��Όc��QކJ7$?��6��jő̭-�H��A�b��JL~]��=2̯"�*���){�	'oIn�n����.q�ѨV�`Ų�
x? u��'�lǤ�!��yo�hW����W+��36���3�Cڸ�&�q��|�U6��R��~������F\���X����wv��W���i����Ţy�N�o�9���cI������s���!.z�f����r�]<��@����ͬ5&�{L�U�Q7�.�΁-[�	�C���x��Hx$��7L*�L1�@d$t&����qj:�l�T3o���wA�i���{�8t�8�X�{��Z&D�{]]�"�;�p�>��$��=S�%E��T�mO�;�1$�59j2��,R�����A���*��jȧ��`��Dݶ��+���n+�#�p�r�)�Ш��TtK������!j�=��-��5x������z9�>`��=Eg���ʲ����
��/��q�*�X�Ao��6�to�բ�={�|쇤�ٯ��p����X�}H֗�a;1��~ö􁩕��-��Ds��#�V��wy�m�&ԅ'M��%jM��`D.����v�3%qɲ�`�z1F�V������.p]�غ�����Q�Z�[yCAȍm}1���";I�n|XSX�{�[�����bKt����&O��^�����ח��Z�H�5!-�[pܚϟ�n���+Z5s��"�E�$�*?�]
�{bq$���]Ȝ�����R^�Q!�N�����;q_�y��c\��{�羗Q��	|Q5� �::^9(�m����^���^�&HY�jr���� �+�Y?7�QX�[�\a�	�+! E���3�oc�._�Ǚ �d���̹��h~���1�\<��]��7��.��3 s�ᙉ�
��X�]aΆ{[�h2��0y�O��O��烂�[Y����J0sc��$e�\_� "���ݯK�̉
R��e�ݩc���(��~����u	4�B1`&_��6.���rù���������(e�[N&_ľ�i�}�Ι�R���9�VׅW;)O�|eS����y:��� ��Jyp2R$
��C�l�բ�,��)<�*7t��	0��c��{|���q�>�v���x5���҈~ׯs&	5%:f�1���������#��lwȹ]_s<^e�.�{���喝":�+g���r�E�O��V���'4!uX���}�朼1Wf&W�tH"R4��ͭnyѹ�6��?$W��J;����L��')�(����S!��O�ε�e�T�
J�����*�53�����������v4���H 77�H�ا&��i� �屡�VI[��j�>�h9(�IR�F�V u��C�I��_o&��^0"!�KB���RT�\5>UrM��o����r;C�����_�H]%rB�o��a�ጰ�����&�SD���)��`u��e�V���p���᫇a�6NU��.i7�B,ft�D�YB �
�'-P��s�	;�Qn�(�˚ FkRU���D��]#\��0��|a��ö����:�T*/�3�u��GXt�D�Q���b8�9\ԝ��'<sٲ��������zv�S��^�e%p�(�[���m,����Lf�d�[��г��Vdc5t���&88(^��{My7��K	F�1� ?6=us�skQ��\I�#Y�Lp>j�{�J_��+w�ᬟ�&��>��~��0�}��k�⛰CFm�C���_���謑��0?h-�B��n`L��p�.i˕�X0� _`�?�L��U�,�/#���J�¶�t��p)R$�u
��}��#�D�f����|BV�Y�I�I��F���i�w���TY��]���_zl����tbnWt�AVqɵE�v�{��3������W�b�TH[��,�u �22���)�d\7YR���8k;!W�H���VX{1��t���y~?GT.��}�x٣7�FOH���Ç�ϳ��h�3���R�^���ﮧ�C��	�wStc����-�"d���ˢ���Ѽ��p?}��P��D�k��ȷ]��͟�]S�	�㈂� �K7�$���>Ť�c�DI|Z��D�V6��L�aH"Y�F��(�B��,�p�>a�©M*�g0���9��匊c��o^�@�����dG,M�k+M8�������*�[��R� ��8����(��A�u7Pqv��%4�,OL��� W�� .�{�r��T��H{p�w��!��H�W%��C�j�;3�U�攂���1aծb0�bb����?�6�E��2�n
�L�s�m�ߙ��6��hqU�y��eJU/;l0�L�ݨ�j����˰�C�o��ϬF���i7�W�Z=���t.���t�F���\�5�z��V�t�Q�.+PʿT>�3��m��Db����^<�/��u�{o�r݂�É��c53�|����ƕ_�-Էt��	�K��������������ʧ�E��M<2�⸱�\i^P"q� b!`���1c�`̹�e�lGK�ƮS�r>�����ې�R�i<W@��2l���!�h R��pk_>�K�4rQ{,:ۤ����*^���U���^��Ugg=9l�l�7��ש���-m����>i�|�qZ��H�22Q.�^t$`(��2tm$��q�^�A!�K����)�]�V7�r�����	g&_!vx���z�k���B�H�eI9ĬAK֌p�٭�2���I�.f|�(�{���c{��]$�Ԯ��3\BYZD����̉�V�0E�or���z���.�AG��+W��M��+IqbY����+���b}��L)骱���Y�	�Tލ�F���&�>�~D���,�5�`� ���tl�M>�r�[���aU�]�ǁq��֐��mc�o��8��gJٿ�Ԟ�5��k+w2(C5����j��$�&k�q����!gY�2����#tCh�pP�I�Y�M>�����Sr�~��Z>��k��Q���$_~\"��s]��O��&"p�U�)�.ӎ�t��adw!,G�S��j��i�Sr˪Ȑk��I�i�U�# �~j;TwC}������Q�Oo���x��J��q�V�m�u�1�=���>ً*��ۧ�A������O��_0�Z�Ď&é[C��.�{���46>����b췕f�N[}�>� =��
EMOf�K}M�2u�P��D8�Oٙ�d�Mh��]ol�y�M���9�<n�����:��~8tԤ�_�4#������٦O���o[���{�,��x���r�����e��֢���%��N?�b�B��q<<�Ti�������"�ن�Q��fM}{��\���D��k�{K�J9wrs��5�}m
R.4S��s���f��C�"��Q�N�S����m�\���*;2��ET` �=�Е������7��Cy�������U���G?���+�(��I\>�>}e�y3S�s�e���
(T���Τ�������!����_�O�"K�AHbX�i����z�� ��]��z�3���G��$�-x��r�$3������H)�H����n���6�Ӑ������z�4.�]���U�����n����r� ��=�9e�عթ�L�D�{3鎅X�L%
�ck�!�I4h`�[͗@t��Mz]�5����'���x~`}G����E�=T�q�AL­d���M�.=��v�F>wЀ�*옻��M��R��~�sN{ܘ�d�LCr�Gh����'��Y?��nm��IZbj�+4}��M.�.u�����a�O�,�tN��d{S�	�����F~/dh1�*��c�{��+���R�e��diw��vb�z�:�(ޞ���db-�,�lÕ�D��2��75���-j������}����	�T�9���T��J� h�A��ls7��x/�$���,�X#�`ei����Eߤ�J�9<gP�)��j�r�$�F��jL/=�(��p�'��bz����x�t'��T�G���R4�j[1��)�$���c]:��LU�TǷ;@.�I��k�%�$�=sZԂ�;�	�X�*�w�a�����f��w��@����`�Ủ�_��x�"1l��q?�"� 1Q��}`qwT�I϶
�n���/�̙[��5���'S��ە&~��3��u[3��d�Z)pU^'
� 4�G,j���D]&֏��ި⮶v>
4ed�nN�6
&y��s�B�1�R��5�$��X�x��y��R\��:�fLr�|5n������l۲�Э��1�y�S�|�5�b]!��W�Y���zѿ��0G���؞��cz���w5f�.1�3|��H��PNV>Wg�:�%c9�ܭ��+"T�.�A_����w�A��U���mib����p qA��|7��d2��a��=����n����@�dK���@�N��I>���Cҙ)ȾS��m�������p����'sQ+�O��.��Xi�␔'��)>�p2�xg��e����+l��w���kDJ����je�qݻ/���k���{�!�!k�۱�Nc��Y\ygw�y���1^�X�^��ɂh�(*�t-�Uk���=YV6������� �/S�S���e�p�7>s�D�t>�ۧ/!Z0�[�9~ʁ�C��|�Uf�A�-�~	��K,�@\���H}�D+�C#��an��u���:>ka���3�7�����`qό&{��t����',�3v��1T6ߠΟ�yK����|�b�wj,�� X*�M��l#$�;���M[ҧ�ّ6�x��b�3g�'�෺��yn�Vd�{�~oͨ����/�,,����.R緯�؈���o��-t�]�a���L��O�,�.o�Z ���E�vV�n�����X���}Q��B��1�+�u��5����?��6�Y�ԫ ��9CI��{ZEi�5��@}Nz� u�,T���@%>in#5�^gŊ���3�@��ү�:�}��ؘ�E��<�,41n�<DF���`�[��p��9:�Y+�G�r����7YC��/���}�Kt{��eԟ����/�UU$aI�ef�z��x�a��Tj�ٻN���W�k�۳S���]�WB��Ri�7x�Y6�_٘M��+�;?�sre׾U �Y�;\~N�4���Bv�g�6@c�����^r�B�"RMl	H�z���$��uL�H��V�o��x�Pݔ�K���������B^�t����2�)1j%ί� ��qX����Te �����~E>�]\ٛ����L�H�E�(�Z��N���zQ�m�=�J�Ȟ���:����[\��0����(���G���U����b�̬�6��d!���޽y<Z���O���t/�(f�<�hS��Λ��0�f���n�����w�hk�>&hk����Wy;O�SHGe7.����QLAD����1��-�zɧM�sW��f�aA�7@���W�#u�t��)���I�	�jJTV����]��`�g1�����_&��M2T��M�&�5\?$kzmg	��/i��F��!�VSal��������ϓ��x{?]�m��K�"����|y����B8��O���lv_2y���cGW��G�d� ��	�{1$,>��a�q�N���-r�����T(�ɪ�!�co��×�^3H��e�J����|�xM\}a�\���ުTk�:��81j5�O�wd�X�}0oSi��z�`�����s����W��I?$
���s�?$9[�%"��;�w�,Q ���%��2��`UA�Dӗ2�2�k�X�g��ٯ�E�?I4V�e��|�u�����g�%�rv+
l&�=N����g����T��h0���W�umh�Fbť�Z�bx�A�J&BL_xQ�U�>�U����3���%#�/�2٪L�9�`�̎w��n�����+�*�	s�W�m>|���M�Ƿ��,Z\�XRL�-�3�$�9����G����Q��2*O�a���vv^ׇ�0�\"�3��;Yq6hT�}SZ�	%��Ԗ�Y���^�,$3"�=�u��z�d-�U���?#�Ysy�]R)�s�f�Y2ž�z'5Y�����������F�?�`�k��lk8J�ϻ���%��e���V>�>�YfW,�V�x��C�Q�z��!*��Bj�L
�� �������Xˢ[�� ���rv��V,"T��0M�X܌�c�63c�aQ_�u�>�uk�r�����9� Rk��F���f�>M�ź����C�䞥��n��U���ʲ��PڷH��"΋�i��*j�^�o��i����EZ���ɿϳ���`i�m�� ���@`�@�$��,5��y�����.J�F��x��F��OԚ*���qK���(�j@AmЈ��x�pL�x�mNt�������l���X]����X��m� �`��.-�<Ҿ��'"r��5�=��y7��N�w�V��枘�����*僦&Jds��b}���:�
uZ�Ґ��1�ul�+S3���L�	��	g�L�?X��*!��y����m��zwʑ�^:"a�A�K%3ny@{�DW+����EO���c� H$�
 ��0Ϻ	p���8�X��N�J�  �<5cf`���U6���0��w �b����9�dF�F��IIX�;���8d�$TrM���e1~�3����5Ie�]�aٯڏ�L�>��oFM;7ΝA�6�;�ތ$[�(���F2:?BW���OPw����%r��,�I��| _��W*Q -X��m�'a��ٕx ��ߙ���{�p��%$�^�7�>�W0����O�PՏ���%j�z�Wi,&���N�0��\�_<Q{�V�KWX�7c���*:����'�|�������/�J�́�)��i�+MKa�9�R�ax�����|m*�m���ܧ!�����V��l�����E�� ��������)ľ�Ǹ�(|28�8�it�C�7������>�)j���)	,i�*6
'�����ZG$�;�!�&:W�|�b� ���[�FAAn:㚃�����NLG'�*����H�� J2��⨊��64_e�y�پ�xF͔a��p�<�u��)���ئ�l�.VkgbV��R��}垱�h;���br���j/�.�K!O����� x�S�+Q�h#�a��X�oו^�0
�Fj<�ƍ/��]+��qr:�᥯$q�����t#�[XdDv\0�]W�D6Q�ffym$OF�?p���#�tL_G�:mYs:}���h��}J�:��](M���%^Z��v;����:4���F��\� �~<��}\���3#�,����#�M����9�n�%ŰE��E����P���v�5����Ǘ�Ը��(�Z8"���V����1|�=���&� ��!�,�@b��ĩ�)����j�s�|8�|4!0����p�J�E���C�5z^ !�0H|�?�sk[��!�UDL,�Ø�E��:�ȖՂ+`���!>�$'5@�YJB��y-vE�(�>0�W�H /�P�w�s������Sy��6��7����e Ż�nk#�Dl���v�'�n�v�7v�<�����@~��^���]��Z�a������/b�$�����G��e1K	�Mb�+�b���V��	^��}O:-g6PbIU�'��5i�������S�ƭ�I83mg�}?��`nRi���A p��_���b� �Q�-Uf�K�IƷR��s�De���D�&2��w_Q����1��3�l/�]-S����LSG�:{>�Zޭ}6K�v�D|~#��\�.����ƅ�#�#�M�����r� T��b!��ЯqKn?S�һ�4�j�s��y����e�R��_X�����������PC'�^�>�Z���mG�=p�T}߹ʣ�r�7�˱�nz���v}@���46[؜o]n����߂1�u�6{�X�[�WC�	������w�D5���	�}�Y1)^�m,��	M�����$���񙌤���Ms���ʗ'0�{�i���9Һ@�n�sEM'J��`�V�1"H�~ľ�A�&p�vד���V��e�FK\i0��|�Y�M>_����-GO��ĝ����t�)��7B�]��f��mƖSq��yS����v����KVr�����u����L�r<�%�F��<�[s�٤��ˈ�����*os�݉���Q-z�r�i\wp�yl�	[0�B�HTP��/��%z3�t2Xҗg��p�3�+�W<�⤴��S��&f݆�w�f"�n���N[u��g��_L�H4�/H���"6�=.}mCDPn."��,P��P�ׇ�<���[��_���.wعA��C�u�+��}NH3�;.2�<(ڦ����h�˒?���?7'��o/ E��kR��܄W0n:�p�ð�e�P�B� ���Zg��E ��ަ��t<Ҥ�R��k� ��].�W��E�O-ѳ�M���ϙ�Q��qv��9�(y�� �%kv�r��2%��EUy`2�����5�ݗj�J�w9v���3%��3�[|k�zZ��,{t2L�}2��a0�)'?����=aC85�ҙ�qD�sIߠ���/@׬_�=柈¸g�4"GC7�����|����ޝ���D^��$J��,V�E���.�S~���X��� /S����Ч�h�\�H'��d�o9l笔5B/���¿̐-�lqEi�˟W"V~�"IJ�'N�9.3�B�8��4��Y��3�Hbۻ��X�u���	�'?Rv�ʡ�3T�E����VPI$�14�]��݄�Ao5�A�F�A�a�6��u��[+��?���N������g}̄��(+��O��	T�*eV`o��0����
�-</�7b1d����J���_�da���[/�0�}��<T@鈌e�gL�L3�(���JSv �H�hҒ��U�O�Z/�_x��|�����$?^��ހrL�����a^_Z�����/qhJ�a�i��a�X��Ts�f�y���� ɖkX�T@2�T�
������w�^C���dCT"yD`�~J���--"��N�6� �n7
z	��D�44����^�<�$��v
�x�_��)�"���ٯU�{ե�t}��X}��	�G�BL�P&���S1�;O��)
�X�s��!�<�Tx���6����s!�!��i��oΫ���*c�U=N��uz����I����k+-�tEm��T����sY��_����%ʦ"���낲pd�?�ͨ�{�U�T�����G�D$�(�c=�F�\��A�
���H������dݼA���lħrW���`l����s��E�1��k&A�6<*TlM#�O��գ��f��S�*�;�P�36�朄��o��B<�Qf���z�Ab�!L�z�gwjf�Qw�
Q@Aϥ��e��BH2��ׅ <������"֏��4Sa�Z������A�D�Ŗ�:i0�q_+5*��p9��"�"m�bޛ���D$�Ɉ�oZƐe�� ��T�_G��N.�
m�%F7���\+ۥ���Y�L�(���&Kp��XV����!<p��ֶ�
1r�������8������"$�Ą�����d^��-mڼ�hC��B���%ē��H�e���_V��?�@��t~)t�IU�)bFY�t�E�~�^�Dy�S������o	�4���<ru���ˍMb[/�%���ߑ_���߫�����74yz��INӅ��~it�rr�DÐ(�cb��C�X�ݒ,W�~���s< j��ǲ�CD0��?$����`��(�7�t�H��G�`A:�UI����1�#����u��>��q ���D,�,�RC#J�`�'�wS���"�w��ؓq-�=.�����SH�l�܍,Y��F�%-fb�*o +�0<�v��tZX�T��^�r�	�İ�[x���޾w7�:�����YFB�a� �\�?P��>���i��+L���Q���;^�Q<�p���:$���TF�f��E�(n���6@��D&,Y</v�>�{9�uh��zq
΢��wL��Qݸs�@����Z�0$e��`'fzn��W��<w3�I:�������U��\�g�kS���-v8�F<b�t&Z�����:7=�g�kT�\�������DP<`]}�a�	4�8�8l��T��Q�}�ݏ���mlQZ��'O�oyC6�:y<��$���#�)��|�f���%vt�+�X�sƮ�>�o�%��#e�}Ь�lH���x��@��L!:n��f�pn�3h�:����c�a�5�������fo�[��1=����LU@d�{�����������2ҌS��A��N5d=Ǒ�~�����Ǹ%���#�M�b͊?�o4��LH����!�V}�� �<{h�__��e��^y�a��
�	������I���L�y�ulh�aL���,B��3C��),r��J�v쟩G5Z8���x78����z*o:� h#�H<�y�NEh#�S]�7�/�\�;>����ٚ_�r�{OM�Q��HR�w�KU2OZ]�!��Q!�r�� n�H�ޕ�H-<�N�1z������k�t�!�����@8�"]�����Ĕ�!y���%����sc��1�����{�C��X�g8���c'�Q=ԜUi�U�pYS���.�O�Y�E͏�S
�D���9��!|��u��<v�������Z�+y����4�:@���z$�\����=�FvhgH�6c��&v�w��'=���>�x�+����sƙA��	G�x>����{��ī���mӄ�/A<�aQ&E�=���s��)�%{Q.���a3�J���7w�H�O�S7���ǔ>5�.�-Q%3@��Xw��x
r�ؗ�!Q�ֈ)�p�B�YϔA@�/p7L���3���^�c��3Κ��͓�딘����-�bO�~��4K��y�_)��C}��Ғ�����A�|�8tY��e�1�At��V�i��r��hT��;U�V�~����H�lq��!�6F���`�
m�LP$�+�b�'T�D����
D����V�rj�\��8:�crA�JaR���VȫƮ '��K�y_���~�T��j��n���L/ �L���֓NY�W8��P��2�t���)�>�����" 5���U�6���'�����r�0�bT�3w�;ʵ�^T�G���p��fٚ~��W�r���� �(m�s�
�S�n��M�c/!5%����	'�5����AS�|u#�ǹ��,WLD�4�{��Q��Ҧ;���M���gY�����n�r���raɽ:D�?��3��/8�4�-B�X9c�.�v���#�<�e��x*+H.B ��#(����7h�����<����C��ځ�����L\�@�qKk֘[���W|��=��#4�Z�hlk���c�u-{b�����7�<�?���NI�*d�Y.� ��%���f,�:�T�_�+@��D���E��T����z�, �.�,a��}>�c�R_���*����p�~���Gjj;d�2y6�|SA���7�e¡8v/F�zEf(^�.����t�d������1���Ʃ��p�X��E �$�lC�΅mx���:>��Lܭ�+�d+yWh��U��eFp~K|ĦMIYc��W���ѳ�S��w;�U�wV[f���pg��������Uc�����M\x�y� #!�]�v,��(qy���8�i���3P[^m�Z\��*��������;J����D&�]�6D�1��J�{P+Q)����a�l��e)Pp�R$�>${�_�h��"�S���/��/M�<��ҹo��_�y5�W#x��%�9qq�c)�AN���M6�P`��L)�r��Vc�I������l��;%�޲���$a�(Y���1,H�1~��?��P�e8�rɔ�&mW =��"�r_�-�@��u�S6����_]�R������Oy'�C��{����J���2�^0'�8���H�cޓ��=���������%IM�G���,���Q��L�4���6����W���?��?������Ω��Z��!Нk>�w]i���ٷ�;{�ߓi�뇞0w����"�~���9��.�KR`A�����C��
�`��S����:��M{�9*�Q3\���+�y+3�i�f���}��J-D�i�^~����i�������w� =��;lx6c�G��g;fU�� cP֩�S5#O�<H)���A|8"�hEirA��}����8,��Y%AB�E�_@3??�a�h-4 7�I��\1��V<_���)7�lN�o{pDZ���v:yľ0������ΰb�)\ֵ�l`xbl��� ��.�O��n��q) u�T�ߝt/�3�|��*�e_�_�F��Cpx"A���HL��4{f&����t]q�6�7��_��h�$Cw�SX�ռ;��Ը}��cy0�����?\�Fi������OBzS�c���m��䕘ír��VR��B��a�JA�z�̳��?N��3���]�c�-�13�:>����D�D����m���t99?L�H�
�Ji�n[���E�
q��}��U���X�s�O�P��v7LE'��������e3�=��u��+?���l�*����[Ϻ����Ơ�7�~̪�x�Z����0g�)o�����gK�����$�Ѵw�N�߻�"nXc��2ЕS�0�=2�!<&(���b���1���%��D��z-��XXl_��؋0f��o]��f��ǁ��J�mo������zV�g���F�c����nx �_����'��U�Yvp��V0�W�8m��c��\j��O({y�;r�.��##d덓ZKȯ�(u�t�m�$k�"Z��Q����n�4���-g�H �����wZ{>J�"g��+��0�)6X�}@�b|C��%�˓�b�O�C�������4e����w�Q��a�v��R�(Lk�9�f�q��\K� {���W�t��3���n��k����ai=�s��v؛ǽ��X�����4]�F����s.Q��nwG3��og�J�j�OGR[,HQ`X㎞��e)�8��B5o���2�ʍN���dY��������}AD}U(AS�D*�M霉X�~H6�ĩdl�P��.����8����"���R��\�p�f-�4ad���^mд��v��l�qbE�:.~rP�����_�	�E�~sI��u��T�SY�rD���
/�v� �R�Tޫ�ÿa0���-���P���/n�\����#���c�VtM���%�a�T*l?6̞��s��[a~����F�t%�<���2E@:��H�F�X�α'�^�`f�Z8V�Xh�)iB7l&�,�
����`��Y������c�;۽]�fjۜ��.����H�J�`
�G����%�&�,IbU��xyS����像G2�Z�QR�SJ/D�9��&��� E��x��G��A!m�;�O���$�1޸��0�.��j�,���"���4h���Mqb�Is��X���A�0�A��3����v�Ţ��2��:�6�z6pc��!�TyC�扽k?�D��,W�����J֟5Q�>'�#1o��n��r��O�rVi�(<^�����׀�GPV�<�=�z!/��`,��%𢶦�9F�	J�4���jt��tߕ]�:8֧ �Z�_K�m~�g��`�3�`�W��NF~���r��z�Au����S'k��e ��$_9�0\�ڼ�Q:����;kه������,G�y���h-;6^�2Ͱ�LA>�l)kA��g8�S�$cK$g��ǘ�;D.�f�y���p]�9:����������-��ǸYH`[�G�*��%��t�UWa5���V����+ƕD3��v�=g�)����(�/,'������õ�.<kT F�����\9T��H;��Q����N��-��xR�N�{ �%��>�bN㺯=��9T�)��+jS*���A>WVB� V������ԥ��Z[/�NR
�����<6%�u8d~�Oɭ5u����
�N�m�]��~\���&X.@S�4�F����A�b���'��[Ai�HQA��3�����y/�#��u���!��r4QȊ�X��d�-�\�q �X ����`�|�A��o1�w����K������}��c�[�2�.� s��F-i:��$I��%�p2����>�����&-��>���_s�4��v�q�vH�o��.͏�����02(�$#4�ABlL\����7���?|��1�%��?��Z4��@�����?(����ٚڊ�Raw��+�A����b	S�m�ﺀ��-WyW���TH!��ʼW��e���rQE
*^��oF(D�RX'
{�gq?�&��S��!oǞ��,;��,�rς!P�fə�I�c���-}�m�5zv��՗FYiΣ%,��y��sMK�g3�u��վ�T��Z�p��:��\
&��&���O"�W�r���,�]�;����J�ln:�!9o���4����7�W�1)��������|������&��X���"�V�*�VʷCq��;��1���?��ߢ��� ��i���Z�[?�f�!��
���7���5�.���rg��vY�ՔNRs�\�k��[�ڔ
KJrV��ե�ld�T/*FD�=�\hD*P����bc��W�g�p��(�0�ɪs4Wu�m�>��y�|5r*�"{W�Փ��h�P²+���QW�;I�����N��F�ǡa���ߍ7r?e%1��f���
��W��y#Y��F��R7Fv�W
Q��w8d���E�҄hEӊ�A���ʯ;����_����>�=ObY�TY�Z�ka
�2�4���q��H�*E��1�/�����ٜʠ��0�j��$ݑ�I?q�L�1�s�n7���1+ I�j��%�j-������6�S!x��Aل�B���J��o�;��3�Q��b~b�Ȗ��"��t%H�7ؠ��g	�B��ࡵ�J��i:�é>����d�d���E��8�=3���-,�i�����v���N�������X'B��ݐ~>�������P�|�><���U�	�M�7��Y�W����:�
�l&�_@�u���~��T�dI�2�U�@b$Q�q|�uDZwt$�Wvڵ9��A�_W6����ӌ��f�FAG9S=�rXp���Uz�<��,0���W����&��Z�I|"��i�#$�I��~�Dt�� �[-
t�����h��qAFb�������hx��c���h��bq�ch���YO�-����>�ֹ�I`.��n�ئ�\��#{�+��"�:�:j�f7MV0���~���θ\�Z� ��~b!��Ʌ�cF����|qʚ'�5�mC���-Z���"8J�B��ʻ�ׂ�+?4;����3Vw;ZF&7}^�ȁ�K�$H�I�����UЏ�	-7E��H{���(ƜICAr.v��U<�U�2i���*�	�(���~�'R��������"w������ԷGS=}0�y�uBC�h��5`��U^'Q�<l�(���ڙ�p��FC�d`��𥡑�%`��Ҍ9����$:C���sh��1*��s�S26ܖ��mb$�O��؝W�����7��I�c�D�:_3��U�K�"�V���Q�����n+wE�}���
�$���$`_��&��'��OQ5�-9G3"z��G�P�F��0����r��}P�^7X��^��%�V4Vx�F������wTiV8g����V��5o�u��j��*Z�"�Mݫ� y�w��t)�
bĠj!c���qt0��0�~}a�465���q��g]��\z∆	\�\�95�k��ȡ��!�Xsl7��.% ^&���nӎ3��fT�yN������@��+�|-]�s�y�?*
�@u����dQ%��'eЂ���|�Y��>�X��S�Q�����
�6��������Ϝhɇz��=��Ȁ;P�=n���������"aW4=}%`�[g��c{�������o�Sٝ.��=��E���p�V?��	1oa6Ph��(������|pBi�k��#"��"�V<Lr1,_�7�B�ә��E���,���.bW	-')�L���W�`ᰞB��=/Ǵȫ2ؠp��ŵ�N���5����˂!��d�/X� �*����HSm��U�ͲmhM 3Γ��aE�ܱ)��?�$^�HO�&���XE�+��7��{��={�ɧD>�%8t�7�ь�/�!zm͌O��4�� 4Ϥ#��l�X&�0^ZS&i���8�<�ﴠ��G2�����$ί��'��FQ.����5�W+ag��Y����;�)���nR��]��3��������D���ԥ�I]u��w�L������и
�=�)	�Ҷ[@��6��N�@LS�����Y�i��v2�XQ���5�=�:(��E�k���"�U[��x�a�p�ȥHу�p%�}����3>�M�?<��$�d�e*�@��\�?T��XnE���ա�P� m󧔌�+��Q�t�OIƹӗj�V�u�̕d�R�q��_yiR`|���.��V���3vW�8���i@�Mc�$(��/�Z^Y���ofUQ22���B����--L���� ��\�Uw!���"w<W"�լ�S�t~R� ��(�e�.y��L���#�����N�p�Q���v��^�k4����� Z��ZG��"���എEr��6��4����zv��S������h*��}V��a���XQ�1�qF�7YoMp��:��$)�/^�Cƚ��m@��_Ż{+ 5���P��dޱ9"�P�!ۍ���]�ܫI�%�,,���js���E��T�y�J�*<EY�M�?dL�%�Ď��0 �S��O���BZ�,V�Ʃ흟Ĵ�(�T�YP��(*��\cV��0�w���J��1�֨F_1)�>Q���TM(��m�5�f���6�=_@�8�ِ�,��B)%����FSS�9�qV�6A�Y>~��oC��l�t։0�a�Q]�n�Ӭ܁bSp��|��Ri4hWS�Ճ<�%���N=��4��^>9�Ю�QL ,ꚴj@�ۋ�v;�
�QkD�	�U��Tg���8NP���
BGD6+a @:��	��JN����!�o� �j*�9�@��o���#���ۓ�$S#8T���� v�2h��핪I��z	[%�m[13)��o�&�E���"��0E*`vH��&ss�+0Wd�p��� K�.�Þ���X�ȫ,h�Z��^y�p��C�z�u�y�~�smm���b18��m��k��8�{9�b�xυ����F7;7��u�\��\�v��e��cś)`k+��f�+��x1"���d�ҥ�(�3��dwE_f�*%�50`1Ht�A��;�i��=��v��u���߶{�ψH��C����i���_ɋ��(��Rq0�)nUH���~)8���)���{��������p�q�*��`W�,�Y��8�����3jί,E��a!ܚ2_�f�f���󴪻�r%�v5
4��g��/q�t<��,{���l�u�{Ҙt��1z���ҙABn5|yk貑�W鳬	�pͪ!;d�+��,%��5��'clA���@P����^`�Q����B Fx�2��8ٗ�z��\��:��,T ��CL�\m� f�R�i�c'�l��D�v���V���K�R�(��J�����goݎ�
��ڳRi0�͟�,��~F鶙S�.S��Y"����~gHG�mPoH�$�9"�5F�
n�0q,*���PJ��x��X�w�yu@�<�����Ve���E ���d7�+�ޫ&�`2�Z⏹i�a�S�V7�R���{���qD��2���~#grpf	��+�.2z�E�A�5t_�wLm�:�4@n$���m@�W��N"�"RX�.n�7��05G�߁O빛���su���l��P[��������f�Rk���]3�&1GF�����|:�~�^�Hg�
C����Ќ9��f~�a�e�X�� �J���M]~(7Qo�E���c�u ���j�����ɰ�����H�o��*,mr=\(�j4D�ږ~�'�܁������c�/���|�cr{	j�w�ⶕ��u)����M�c����ǜ���|";�y���fJ~՛F,��5'T{ROx�x��]�*���'"�S��F��,��EuI�!�]r��N0U}<�ઐU��Թ-7X�gk�QވڟcĚ����s�ϫ9��VkA
X�5����%RI�߄�O������} {k���惊-[�7�R�����BtuC��4��Lr����}�D�B~���⊾ʓ�����S�d��e:�0q�^�vu���Ii�A�.?���To�&*lqx���j	o	j웾�;?���������F2���r l�T��X���9�4Y�΃�.�@gg��$_�7H6��\.,�e��ex��s�P��)�����R��}�߯�(���?j�:�+4CT��0�m�*�I�o�ũ�O!�LDQ����0K4H���#vtl�$ϥ��͝�{jnS�Bm��l�.	D�\���F@6,�"`f�/sϯ�Rǡ����	��p�p���"KK�x��0�P�+o���yD�:����S�Ė��3ǋP��P�Ŏϝ{g��D1HP6WCB�+���j?G�0I�|��h���k2��֬ +���h�*G�;ҁJl��
�$�/S�l��a��{�B�;+ж�;{��%nS��� >�L����^�X2��N�;��ھ��z��K�9N�>.��ʛs6��{;���6#�*���8Z;]}�J$���cN��v��*��,0J
��I���UU@�4Y��jĻ�c���G��V�@�<TN(|�>C%3�,���{�����k__����`����ف��My%<��M-oR���"u0�.�z��_����QHgr��k���r�Y~ #7��5W:/H=y�J�#�%XL�Y�b+z��c�:����/4�M�wk�f~�t��i7գ�=�R�t#;s
�qM��2Rp]\��?����3�UwE�]vF�>������v��ZK�p8�?T�"��M�f�`���ð�wsz�h��ܛw��V�ϓ������W�l�I�Y���XƐ)�	s�G+�3���`>�i������Q��<+e�ʣ.�B� jb�\�`���_����� �A7��9z�8�3��ϊ������Ȋj����Nu��_��}�_&�.	ʳ5cϱ�g6E��q?��s<����B�8.�;��O�6�`k��M��-p'����l	��O�넾&č��,b�$=	6��{+�x�,��FBF]�(lڑaXӂ9�Ȭ�^+�%����͙�^Y��F���u��rbլ7L3�!lH�o~^���4s�M�1�&�����pS�lb��akE�Mnl��A����SsȦ�[�廉�ӥ<�Ĵ`ј��f��Pe���.�����u��M%w�)�xy�qG�n�:�a��=Rx����ܪ+7I���87����-�p_�k0�{$����1���r�D������ڄPm���F>���~�L1A#��G����%�8]�4p�Z��Hʄw1`�7�\BHo
&U(ђ����L
.08��?L�>���b��D�] ������+��u4j�����	؆+R�K{�J#� �Ԕ�������?*|C�~s���)�Yy��ەG���Xc��-)Y|1�u
�z/��HK�,�2q4�K*2t�	�N�7�K+׫���><��Sn�ލm�m9��C!;�q���ҰG�u|���ٳ�����H�1&>T'H��y[�(�#��H����3/��2�����P�&���<������l�"�k��0�͜|��N�d")jr�@�E�XT�} uN��'TR�jZ�A޺���|�jǘQ}��-c�Xϲ�J�Z�m��@�ě�?O�Ȍ�ӝ���{~�=h��EHB�R�n�~it��ʓZ������*�>�6A��(KU���Ue�#�w���漬�b�cB�{|j���M�ծq�\l'PNzw������"���^�T<";��V���w���{l<c4���.��W����]�~�2������<[Sl�4�]���w#�/ujّ�ˢ+I��Z��c�X�vT�9əx����T�<)�{E
���:���u��m���A�/߄�l(JہL�;9��d*z*QƯg�ݚ�ަ��$�$��0N ����U�!�>�z���Ḽ��@������A�L�J�H��	�tV����ّ��%�ɾb�-��K�F�(�-߾+7$-}�K���\_Xu�@گ�1�r �W�e������WZ5���ǅ$��aX�s�tR�1ԥ\�'#��E� �V����ȭ�_�6?xJ+�_�����;�^}��vs�4�r��4�Fe��ײ^��%.�U'Ow�Y5l�C�?X)u�	�k��MP�=��j�������H��*=��O�MW�\}]���Z���U�ZA���g1�&��@��)�80(6_xګ�ε8�����>Z�i�)1U��^���Ln�b�УL52ޖ��;����3=��W`����:��w���B��hqۻ��}o>6�c�08n�ߎĎ��1yR�f�������J�xIO�۵�U�2���u ø��
̕��D���(�q�
_���q~f��JA�#�k���Bwp��0z8�Z�*N7�C����1`����GP�w%���n�KC<^(0*r���0�7��V*~ƨ�� �?������MfX�rKd��:�����N&��7��4mD��ϧk�2n�<]�A㓖�>m�,���2ӽ6R�B���|��Q[�M�o��q�����x��i̔1�Vd*��]���E�t�L�p�@�� /hr�[y%����5�����
�Z��#M� ���F)H�śD�����0�Um'��1��H*Z۰_��W����WI����9��3��	����ŕ��}=����?�_��w��e��t��V�ޤ�>�lU�Q��\�9�U�;��)�^r����j7�*I[>ʓM<���7e=(n����hv�N�j7�xX ^�@�����®����k�3踢BnG?ť��3�O-a�����{Ʊ}��i[�@Y��B� w�!�-fo̜���x!���Gf�4�"�p�%x�C@ks|D]�ao{�VB޻3�?`�9����s���z�f�`ؤ:��@�パ���(�Zd���{�IHK�擷qsoL�~�5��	6[�U�
�ZNگ�^��H!���հ�-��|b�c��L��Swq�~v�~�#ۂ���(��n_�3�Uݶ�o!�|�S%�[�׷�LՐ�R�aw'jгJ���g��Oш" vr_[�3�N�󡠄��F���	�XW�q�������_w��+i�<��f`�w$�m��L��+^����	^���
筩q��T���%e�%���2�+f��Jz�0=��W�o�=�-Bh����S��M����^U���czX��������H[߷M��;<�C^e	��g�`�#�J������T8���'�2���u�/��GvE"\�*�߃n%����2�N8�	���ƃQƾ�*٭�܂�̌�S����F,8��Vi";�jS��f/f��rLJ�e��>pc�+���x���f�����#"���H�7�+*�a�˩J� ��#qa�G�Cԝ�I�+ ɵ"�H�������j���W����᭲S�����3���@�ƙ�'Jj\N�*v�W>���,3]���afZ�����מ|�E*Q��+Ε��P'�&Ho����F"�Ip"�mʉh�&c<�����/��4�-�@�Ծo�X�co�6��زGA6ȅ�y��@�a2��ˢ*Ǭ��]�Y�O#z �<xV��u*6(7r���q]!���8{�h���0�����(ӛpXU�q�U�(gD�@"�}���]�4ko��~"Z�{b��&v��Zr��U֪BL��t�-�yc���U�Zb���F�˄#�~����Ѡ�I��[:'�kB�+
�-@�Ƌ̏�����+@L�U^Ix��7��`US�l��D�{�4/ָm�3���zO��;]G�٠�Zfp�e9T�f�!�ee�&_��Rָ4�.c�s��(���4i?S��ݖ�+l�*k���a������b�BzN��9��O_�vQӤ���}��E*ŵ�kw�5}RϚPv%X�(���#ޜ�5Ȋ�.#�D�ɔ�2���%	��G��CY�+�2 ���V�`�\���v���v`Sږ���2Ej�ɥx�1�&I��� �O&D��E"��wx�㊣� ���F�>��܍T|\e�y89>Ǟ�	��ýF�l*2�1@T�.%@���-U����`i�p@�Հ`����V��^z����7���K;C32"���Z�Q�J( �3���{۬o�s; ���*�.���e���&�g�!�&��-�f� Zƒ�ϏB NY�3�dYv���Śs'_��Ɠ�3�/�F�����$M5@��m9�M�̱ �T;�L����?�]ۋ����ۢ��J�(��h��ˑZ�!��w�{%іi�>��z�j��b]-���yA ?�z:�vO�%zW/=��S�@��9�d�����"���.t4N��d폀I�zu��ч�ˢ^H*��I�X�2�I =è�#�S�~�rE�쵸��Y�x�Up�m����f�5b\�/�3�o����x�
Ȼ	v5ig.̘��A�#�Y~j��f��{���C��n���/�C��2@�)�A#���&�����p�=�2=	��IѬ�ZΐK�2��J�����p;�bz�r	Bn8�������ˤ)�_�<ݐ��>f4CE$N�-����1�w�]�GVĢh4^�*�,B��7E�xg��#����G��[��96��:�����XD �����ñ����,��}�����v4���)��$,k6!�J{y��c�7���9:� Σ�\N�'�dA���ik�Wμ~,t`��i�����ڠՀ��|�yR�AP�脵q�;OlI��h��8��d�'asF�Kz#��X�=���&�nد$"��~��+mz����,`e�j��h�Y�� �~b�7��GѪH��Zn���>�2�DV�����,�nL;�)kFz��i���0E��j�L��t�G��#�ug>�8DkeT��G6��,Z�2�kv3�4e(�Kp7���(y�q�s	N�.=J@a�K�L> �N�d�IG��&�{����7s��b~bRٻ>Y�����&.���e~h���Rh0Y�0������]5��gBl�X:"MVo���G��?;'&=��fɬ�XKfd5��NR�zc�]m� r�@Y���dl��US�
��}<�%���\���h��Z�J������	=q����P�F�w]Z@Y��k�dR_����{wF��x�|��i��.Z&o"����tr@�i(�{�x좚(�,v�/}���8X-EQ�s��ɤC�fZ2���nwb�yN/�J
�s�{[}wN¢�`w���֑=�;F=#�\���h�O;�a̳���z#nM�D(o��L��o��\#6 	j�	v�%�:|�S�J�U��k]��0���~w��5�ݭt'�Ի*&�t/(�����;n�ە�ҫT��	"���P��3����џ��.qS8cp�+�H�''|a��=��.͚�`�E��J�G�d�LY�KkC:c�x����k7k��3̗%d�:,���m<_NX��7�(&�S$�,��>pXe��ʶ�Q7+����,����4�C�H5��D�gW��d
5f���z�Cm���Ic���=�I_�&felB)zYGh�>@�+�0
1����N���g_��Q|�4
��Tx#�ˊ�e{�.�=���W�&hB��P�j��߈�B��m��u�8��\�|RGi�������e���>]Q`�#ߥ���,�#��N���=ꃝZM�=���$�B�4�������衜c�rf���@*{�T�Z�8Ғ	x���<�~���_�aߩ�TҺQ;�G�(�I;��+��\휴���T�:걼W���v$����iҕ �~vDچ/�ǦE�3m��Ѣ{�ǣ���>�A@#+�����&�(Q�P�|�޵�+)ai���]����)�vQ�Gf�R��'�l��J�sye��ت�~|��5�KN@��Zӆ��q�}�W��L#)�����ZjS�������WS,�Q��x�h>{���9��05q��rDs0�r�4���_n1s�z���+˟�!�&"�:��2�g�y�af��ߕ>8�x% &��-(XJs���O�Ct�9�%�"P�� k��^]��#��	�&�i�-�%9/F,m��*�t*R׈m�v�+䣶�
P�l�S��C��;��^�e�:̝�b��� ���w��yX^�w�!�~XG]�i���sH�J^C���fS����{�Q�I%!@�Ҡ�F�U��n�JB,N.K��B������nY����;8 "x�?����x<HߋY��L�,�p��>|�k:�����F�^ɶ��#Q��h�W�����ӪM�\�Ndc4a�t�@���,��})0bB^ػ�׭�@��>/�_���گ�x��GOʅɊ�Ry�y�B8�?'Xm��qH�Hy�rZ�����2_:]?� -�ZAx���@�*%p<���%ET�ӪQ}T�����0g*/����0��>:�A�6>� �S�\��/��%�^���NƓ�ա`��;t�w����WKB,٫��#���;��q�����N�q�c?�/�N�Ui� e��������"8�\؆���	!mLx�İ���K6��TN� ��m�����6����8�R����4�G+c{C,ى�N��x��\�Y���I�G�@S����o�����.}yln�B�q�G#��l%<�ĩlټ+�����*���*�Cޑ����g��P`L6�q\('vJ���^qy�x��J6&CܪC�諦2;#�.���m��Db�VB�=IQ�3l���D,�����(��v[�S���6X+��#�3z橭�zg�txn��T��^� m�Gw���z6Y/\�e0��M�%*b��5E8peIl�4��]FF���c|�E �ۈ���\��}R�x�t���,��{�b9�/9@������s� �Sj��M�aݿ+�����6ESa����r����ܶ��Zk*z"��R������� oDPC���u��U�Hli�{��jlC��C���hGK�IY�/h�\'ۇ>GW&E2V�E'IXm�k�x2�n�X��_���84H*OB�F:�+�g@��uԪ�JP�Yy�n��c_?K`�^�s"cC�4��̋��lݝ�h
�H7C �"d�f5���y\]bU,H퇡�t��1�H�AI����(}6fi�����#5��(X���'򳖀����#*��֍�~�[�����.����D�o��vM���@lIb
��\=�9w��u��9
�~*�D���3��ܯ�n���W�'vk��!�2���׿�ن���#2co��])\�4�*iT"�"�Њ$�kR��ֽ4�ͱ��B�̰%?ohfT��̘�����4�<�iM�\y����/�.���ܳ��gm�G{\�e�D�͓��w ΍�L��5��؁6p�y|p6�֦�:3e|lc�2�=�h�<$���Su�|k#X���/ڦ�)h��������P��k"֦4]��������i;py�z�yw���0fG�t'������4��tG��;>�lY��-��A+<���ƅ�2���� s�I�e�i�d��K�/{�?C{�'@U��>Q#80�Ц�'�w���o�͘}k"��7� �~����&�*�4 Hc�acƅx����"�|*���i�W�Zv��ӝ����[5�m(���Ǫ��:��<\��)�<�I����X')�KU&�Loy���T�^������&�C�{�5lzǵU4r���OR�S.j��,�u!�P�ɒDy�V���a-h"��G����i��_�U+�����P_���W�H4�SJ�ŗ�wh�o��aY������S�+���*�Nu���{�����Q��z��mG'L�Ǔס����8>	�\����g�)-����;��H�
��4
2�{t�sµ�F8��+ϊ-"�C�6Ey��\腚:�%�Q�����ś�Q݆6H�d8�N�cV���B�"w�7��������	&�ޔ��j��m�x����;4�m2!���i�'⶚b��.v	`����a��.�+����/���p���\���R���k��z6�@K���ɋG
���"��Q;��q����S�J�J�s w�#���g���8c����`��U_ ����D#} �LmBުظ�eV1a)a ǝ��f�?A����Z��;9)�~�iѧ7��7+'����E�FD�^����S��6�\L�(XM6,g߸����9�+l�(��zjJ�5#������מc���.��v���-f��xjn4�1�˞��~Ɓ]���7�J�$XS�!g���I�nC�n&���@.�ׂ�V�����UQ\�0�G�x���N��d5��}�)���p�?�����'�Y����c)Q��D������)��o�������
)�%�-����ޔ�
F��Q2=?�h�k@5~!�J��V�ԯ�!@՘4/�X�ؘ���QEO����F�]r�㊫`ENg%rW*�i�����|�J;a=����)3���
�q�>���������S�U<_l� �v���b3��ax�
�������s���b<��x`Q�t�}�)}@��,#�k˖���k=V���3�tH��Q?�5��7�߁\Y������3�A��;��|2�AN���O�D�4pS�)��5n����@MZ��F���e�~��	O������(b�u���=	A6�Xc|Jrm6����=�I�΅>��S�*%`4��gBuE�P]�D���Z�j~�����"��k��.���h�p.Q�C�Z��B��DL�s��aqϖ��91�f���Dd��ާ�:�3�9ak����2�V�ŉ׼�:(1B�B<�I�nu���[v���>dx�H�G�%I�ie7M�fo��
E�>Cs��a($�ӛ��0F��ŭ	*z���Ka��.��ۖ�t9���N��(3ŗ��5�e"�i�SV��c��u)m���|�W�K�Wi���e��'G�C���p�4¯gg\S:>��j�s���'�th;�{���M]�2|f5��L�������,ܱ�s,�t����&� �W�����9 �C��p{:ݿ0bouJ=�F�h]
���x��;�I����LB��_�Y:����ė�m�������op�s�r
�ıR�W�Y��!�'�RjЍb�.�^(	D� ַ5�(V���$�����`k�ez�^}?�J?�c�^r�4�,b6އsӃ��Be*#�i����J]��$�uAN���x�R�Ж0��z(����{���T��o)����#rA�pH�K=��i�=�N؇G�A4}&�Ca'<�Q����Y��Yb^�M�A鍚�+��k�D'�r�z�r�r��Q�+V!�o����0��C�R@�����B�km��{�+����4��1C�.sˎY��m��x��i��Ը槡M�V�b�E���{�+z4�}�/�MF�:���<d��{�GKj#�P~Kr�������7�K�5U��y�Z�9� :I�SB|�8&�	�F܉�$�[oO5H�B��6�}�~gn���
��J܈`�֒:��Y}}�o;��
9>�P{u3ъ�	����`���Xר�yj�K�uw����Z7���U@
�C����@e��z�l������b[*Lw^$M�6ω\ahnȫ��΍[T?~}�?�O�I�VQ�Ղ���f����违�	����(�D�ű�k�]Xr��T�S�]�v��K��
������u ���<�4?*p��L�3M��l�Q{K^<��4�ri�[���ɧ����Q�=-�k�I`q����f���qǣ������mmT��O Ct�[,�9��G�������[����y�b*�ݪ��&��R�a���Ŕ%"Sp��٨�g�A��=tp��>�~�Ь9�����x�Z�+O=����&�T���vu��\bmҨ�i�و�F�|:�_A���>P��@�Q��\�s�c�0�]G}���HLc���2�.WbZ��`��/��L���17��O����Mg�5��ƅ�H��ƹ�I���!�U�w���,����9�f���#ht�l��p���S>G���JH���{�Q�)	�^4��<I��+���W���WnA�}��S�S�" �w9�}Z�o������(�<���4(�2)_ؙ[Hխ���.M>�]�[ž�V}*��|%�=}���J��Km��t��d�3=-n �ƴ�/���A��崱Wٶ��Q��l�e�f��#>��s*k:�b;��~%�p�hT#���/+���R���h�ø���.�8�y
�a���_��`�#<7�jwD�بr��a���q�D}l�^H��v�K��Qm�̈́}ޟ�(
�']9G���T�X��[�m�DM�X���?#M�%��\
I��R�f��n�o���D�P���z�#	��3WF�<��Ѻ�1
*�����l"����~"��q� *xdq1�Pu�Kw1����j�_�dm(H�%��F��c+�k��ė,I��$���N���۫A/����CT|C�ٔ;P����g��`�!Ki����Q�4D2z���]kUΙ�{���b���st�Շꇆ�4���A3�Y���F�Q0��}���b�fb����)1s�׸~�^	 ��l��hcS_�qb6*�H��h�P�v69�'ϔb����������"77q�Nr|�x�6��h���M��&���ɽ�N��-΍�/N�UF�rظ���\�l[�-�r)�����>�d��8��+*�}�E����O�ğs�vA�$�ugǋw��RU�qÎ�(hd��h88~�g��:�{�(H��l��_�z`����|�D�8>}�Ά�}n�UGif�pizܝ�A<�
�>���.+���A��������jNPw�J����L~�͊��W^>(����tZ�Z��<O@���͏�DC���9Q��L�(�;b�~��h�q��j��n��7U�p�u?^	���	�ǿ�,[j���z|?#Cpe�v��y���_�d	r�׋2��4R�7Ne.�x�,7�;��Z7�c��� PmLj��*�kP��U:� ��WK��u���9�]�P�H�%�(c̝��}��ox
͒ 1!�K�[�Z��D�h��ի�´u��CR���5!p�iv{��+Q��EB0Ci��YjԳ�l�����`Xg�V�1(�ҢZO.���]��ߏ��iT�_�e�V�l��cO��J��T�"5vM��^����c�/91M��9A�}HoA���� �d��8zOT�I��X�$<�go��xi?0ON0]=�W0tVsW~�dQ�P@n�S��;��gܕ?d�m�i���no}�Î�#L0g�~m��H5E"�l^M��^��EX=ίV�w)��E�����S_�,|y�T%�όw��%�Ȉ)�!p�Xм���%=lU�Y�>�:�[4��%9L���R������#U�>_�v.���ȥR6�������r@�����4��q`"�i�.�" �>;��"F��~K8��o��zp=-�Xo��#z��n��w��,�I.�/��*P`�Nz��h_��59���l�Qg�iǁ��=�¦q6²j�;��qx<�X�;��i�?��N7�\Ї1�h�.��h�&>�``&_zк^(e�h51�5H7\D���u@d�S������u�E	���Ѩ��Fvھ�l�E6�� ������1�����oV�}{?���JT>;�Ǫ\�T��Ky�}7b4]�6��Ҏ�o�-���� e�3�0�rW�݆�?�Dr��Dw��bdI�5�_1���5��Jd�r����'bC>���T��	���7ѲPT�k����\	9����v�	 �ϗ�)��F�F�������@h}����G��:�!����:����� 4�U^�7s�6����v=k�բ���NZՍ�3�90��Fg��ٚ�uDucu��Pn��O���$��]1�:�o����E�R�Au�����Ӎ�z�wg���ŋ��� �	`Y3�����X0W�Yl� �.3^H\�4�B��p6�/�0�;�w	m���Zf2���������� �o��7�!W����C!�~�|zW��v�O���G��K�+��L��H;�Bc�X�Â�
�6���T%�{X���xN#_��"��E�O�0hB�׻���E?IG'p[\�T���߳ �`Fs{��kN�2�ׄ�I��uR8G�B71�gfD����ib�|���������,��3�CF�8a(��杩ܫ��]�Q�vmjJx��{6�B��V��x)��c����,��cn��&j���XL��AHR���F�EQ�M�52q�0ٗkz�sn�=�7�LIZ潍�۲���@��N��7z�ϵ��\�B�;��> �R�z���FcS���<%H~�"���wh�m��X ����Z��o�G�1ױW�-@��������ʍ�	>�m�M�n�����`���d��#�>e��Y*���D�i�3��4y"М/��("��>��jiL�W?��#��J�-�BZ,J���|盀��^}�ڏ0��.�f�I��w�U�\*�ǻ��A��q.�-�OK\р�_�,�2z������6o�Z�q�p����ts��Yb$d�1%W:�|&�`�*y�������F
<�'C��N���a._�q�\��zʝЯ[L�9�Bl�H6�zq�q���|+�Y?��"AW>��������U��C����=}�i���jS�=K{c^����j�؛�g���&c���������Fu&��SL��;��Z��,x1���� �g���w�W��ǝ�8W50�S�;)���&J{��~��V<����(�������4a���("�do�܌��o?�?�Fo����	��I�^V�K��\u�2y��0�ڤ�V��k.�~�����n{iC���~���%Dr*��
�����bH�i�o��]�Q�xH��Yks���9�Efm�}�<��~?�G��Y�� >�U�$�?� �i`������?���䥻=["\2�U���@��I�g��������/v7�q����!K/kh��=����-������o�&O7���C*�������C6xt���{j^�zRa����������D��@��Ș�N�~��d�'C��o)ё�	:R���p4��� ��8/b�B\*�ӣ�h�\���ap$k�O�6D��z��sń7h��ꭕ�(?�1��^�/ǳE�H'D�i�/Y.�pS{�V�Y#�6֙f�S��\q{HZ��&�_�K�����<:R���>;��Ө�������Z5�i���vtf�, ��+���郴���3��+8-��c�yt"�`5�)��D��ۦ�����)������X��w���[}�e ���kW�^�^�ӽj9{{�|�6Ǐ@�����9?n5�U;��)�el7L-��wm�/�&�t�\��y���#�'��Ņ[[TҤ�ޠ��e���[���zj𯭄H�;O�����t��~.���Cq������GU�G������L�"¹��[���W2<�>�����.`��.�>��C)�LQ���DF�,y�Ɓ�H=n��H@ʺ�������+�ҳ�nI)�!?��V��EX��Mj��(T1T��u��T9akC������W+�8f�ܤ����fz�B6��՛��v�2n��ʣ����u�2�h��C��-ZG;�T�3��əf����< ��y���ܟ�ì�,Z����:�2�ͦ��� >���e�9�r���b%Bc�	CQ�>3�۝޶>I�Xs��P3)]M����lb�~�l�&P�H�!1�sja��՛]r�Gܛ�=�l�LW��kV��������إҒ�����8<�
��N�bz�  ����B��ȃ�į��:n1���I� ?��=ē�i��F�Q��=��:5朸.��3�kſ}/(�[���Lu�j���E
E��NCuG�]��9����48'[+z�����;|E��B{��:��4	%23aZC=֋zu�����aЛ�X{vy��`D�Vj��&����Љ�H��6�Ϛ�]��9��X�����U���qX
DdOL�_.�/J�)*VH��u�4!\�D\8 �w+��q�e"�-��2�rB!�����S��0��QBq�����|y\f`bc�<N ǰk�~;�c������-?}�3�(W�W�,:|3L}����̱mu�S�{�F������G��\����M|�BS�%+_e&LkR8l=�U�AΈ�\\��m���d���͎!.�
*$}��@ԃ�T�R����m�Z���2�k�75yT� m�y��:�(.�Fs�{���.��\C��)��,����k���>u��;-����o@�9M?*5h������5:�/�>�������,B雹AК~靏����Y� T��1a�ߧ��F�����U	r��,��}� ����۔և9)���}���;����JQkm�����r4+B�.>�tG�:���UOa����ڙ��^ˆ��1lM��� �JHs'�[�$U���Κ��¦�[� �����c�4(�y#�-�|�����������HhEg������h@$Ӎ�@���W��E{����-W�U�J�����uGݭK,o�.�Fg���NW
�B/h�C�� ���
	/�=EeN<x�W(��
�������8:�+��9���95��~�y�кz���s7�Mf�)c4C�BF!zҽ�6�3B
�7�!1n3u��*a�0k�O���XOBɀ�S.Y�IV-����	5���P��{]jbX*�Z/ ��)g�J�Ǎ����n�k���Q|K���?�9�)O���R%��|5�`ϟ� 8?㖎R��d��^}�ӱϷ����vyU4��~Y�1�Rީ��Z�����d�d��n�O�549�,sSr�l+�^��N�v�a���ʎ��1њ��ԟ'�C��!�}��|�=�2�O]�%���6bKD�{�(;滋
�j�F.12}����'�Q�Use���uT��/�j���
e��,P>�W�"����I�:����/�(c�0&��{"��b6�Gx`�QX�<,�xkh�x{���dA�T<$��7�*�X�l7�tI�����O�q&�a�Z�9�l���	o6���v�:�	_qrh���S��e�>��Hi�����*�p^�����D`\��c�cG�*7�V�����+��!צ�5��*��Km5.�WkS��ԑ����'I�#3��~2K�`䑝�(s"5�4�����$�߯�(^�Y`G�bp/$z	��I�ayV<��Y�P>� �z[��U]�V��n�g*V���[C�<��!
l��F���& �V�̀] ��Ѩ�2IN�l���t��s��▆���%�fM"��������z+�/��u�
���2b�0}5h@X��hI�lo���H���֢�3��i��&��N�*w��'�j}me�����|�[
E��TFU9\b�c�i�
~H�n��0�*�9�[#Vrpij15��;��)֭ ^���� ���N���k0��SZ4|�6
��=Pν��U�k�2G2�6���IB����%�ߦf�z.������i�K���Q�ٲ��5��.�ܓ-��]]:����@�)!WI����ڋ$�P�G���p�}S$�c�v�I�0�Sg1���" K�(����@.c���[�A>p:�=bu����͐.�f�F���"ٷ6ma=����������4)U���1�j��^>c�y:�ǫ��,����#��+�����v��g��V,���ђ*�0�<��	���ħ�vn�0T�I�2��������� �:Xvk�u�/�e��i�����펁�L	��cwO������t�_356��nL2 f3��\�1tf����~�M�Z%�����2�Ӽ�X���[��P}���o�����~�a5�$҉�����#-��֋b��8.l�r0��ƽ��]c�.���V�p'h��͡ʱ��Qǭ[�4~M���4�|��"�����5'�`(�":��槂k�#��y�����:'�u�C4�Ǆ�ik���D��bp�#7�D����f-��&$�:�3��}�άYd��-��sڥ)!G �{�37U�����ל`q!�Y�65n&yu�:k/��=����Qz�����o�iܿz/S��6n}~`�q����I���`�df`�M{i�EM����0��/�Ax�i��C�R������q}�9R3���i��\��W�����2�a��`�'ȘV���-6�������,/�1��z��e���,h�C�y��Q)�*\����
Jb���E׊�&�/���i5�����h��j�?�D�{S.��p��Gx1�u�*	��U�d�<=0�d�)5k�U�P��Y��v{�V�=�'>�8�S����l[�E��������H�o
����m"M<(�u�<�*N1bذ���/z	����hn6�*��?��Aۆ5$�1�7���~\˚T��Ǖ;f��� �U�����l9C6T�d�H%A'������F�����&eV�A�-�؍I�Яe=}:u�-��Xy�^f���hƭ  �ۿ¼Z��Zi�=Gk�h�W���`�S�Z�t�=�u;�A�1я	J�cƺ I�e����0�
[�X�g�m�&�1�>GJ�N`�M{���m��D�&6��w�b��;װ�,�]�,�r��ns{��a�-��?'v'�vT�����?œQ;���1G����!�8Sm>��q�Y�����Z�9�&g����^�ē��QX�4���Y��p���V�[
�u�o'|�k��ݙ>5��ZMq@�Ƒ�B�j��c*�o���V�Aґ��9�k���H��7�Ԥ����ب���E�ӬՊQ���¯��!�,7���t����K�(��Smg�x*�8������i�&d_.L�f�����iNR�������t�l�W*��,��w؛:�<�x��e ����"�vB��Q1	�Qs��Tx|��@U�P�+�9�"�[�D��5��I��{*r�3a<����ə��*X��u�D�&���IgĨ�[�M&ѩ�Oی�?f��X�6�s�n��E7>L�ov:�)��Oa��H��,��&@���VW	��r�z���s=�!ȕ�׭��N�(�����z1�-_�R�d�K��\�����aN��@N�&S���(EzL�)��q�C_���_�&�x0��#Z��O��jXV�<��r��.6�]�1gtۍ�iY/M���A��~{wM�v�I LK	��E����ĝLçq���t���Y2�sH�ȺeT�/�0��O��&̖���#O���^[��\aA��c��&�O �����%$��9L�bLS¦�������WjK�ܷ�o��T4�*�8�E=wJlt�a��(�Q+8�51�0i�؈�a��MA����P5Y��g����p=�/�r��Q�ɖ�>��B+�j@A-�_��0Av�'r7G�q�����_�#���.P��(����8���/��Ү���&�dchs�<F�J\��q9*�Lˠ����Z�ć���c���၅*w�	D��v	�<L��E�Dʏ���ӃtO �j��`o��º	r��9V+0��\��U�Y��r��Ic���ę����츯/��`M.zZ�R�=/�M`	'��6��6�O�$��,(Jn��	0T��(�T��&�WWz	�m�_�s�z���Մ�(�XB����H�x�$�� �� �S�:7��n��_EЏV��>�A�=IE&��#�b3ǰn���_a�K�u6kA���MJC�����HT)\[�3U�>w_���
a��-X��^�C?�}1�v"��V�>A"�#Y<[�xid�,&��Q:~Q���Db�|�;ժ;W�W��ܠtI�S&��BE��EQ��*3U���=��`��:yg�<�����NP�h��eۂ�m��n�/��S�M���?9aH�e�$���X�o�I&eVs\�fq�\��s>��b�,��ZKtiP=UX�Fl��$�gWk$���_�J\5�+n��z�r�jT�`��M�������xu��W�D�Ww�1��w(�.q��T��a	�H=�[]������7O��$����b�]�ޏL�q�),�Cm�t���șow.�8���*`o�v�<��\�[L�E�����8�̍#�࠹��߃ْ��n)ҥ�|����7�g��H�.��lo���[,�H�<P��l����RV2��d$D����9� ��Q����CzǶ0��¢k���J|QWy2ūKWTt�����w���]/YJ ��T
�#w ��eA�ؓkS��mϘp��@�?I�ݨ����It?Z�wK@t�#����v6e��K�t�-Ex�Th$�j߭�.�It�+�����(f��mD��J9�,O���Ů����@f/EZ�6�Ex��,z�Z�¨�
�F'˲�I:�\5����bx����Gt���3,X�����x�����7t[|5�'f{���֦�S3�# � ;Y���0]�F�I{����/�<єB���;��;���q�+��Thz�9S"�F��cƎI�r���9	ɐ���A̕�頪�y��,���By��4S9"�-$}�a9���yw�	�[�Up� *i�g�f�����F{5����E꺴��}��8,��L� &U�.?�l����"_��K<`z���(�ms�	���(���*�g\�*�G(�̵,⍠\�~��iO�(D����Mh�.�E�M�2��G��cb�V�9,���F$Op�]���B�GƇ�$��c��L<�ń���.?m�|�ie�		E�+��M���[��b�&���	|��ih}�w1��H+;�#���Q�P��~��tPr7GkP���^&h<Eo.����W�����*J�i	�4�'1�ݾeg��ң$m���g���@�Zi����4������h�wd�(H=�t��� aymt�r��K��4;���5��n����1�N�q�� �2�2�Wb�p����iZ�?^]NҸ�D���3ӦGº�k�#s��|欱˽�V��^�-�Q�s
� �U�7���8oAݳ����(#e�sc�@��k�VP�Vl�l�RZx�C�o��K�U0�r$ �L7����*�#W>��m��� �S���[�k5+�R��/�2�-My�n� P�5:oQ�ˮ�YP ����T!a*���'lt�vk�f]%������ο����j�^�?=����J��G�9�n��Hѩp�/J�C��̂���93��K�ߟ�x	�M
����J�����_|�H��E�BkG#l�3�w.;�/�e/�%.����i�2��ؠrhn�I,�V���1���V|E�k�+�d����K5��(j� ���� ;(	�����P�h�7X�-�p��/4	�{; �IE��*��0`j���B���8�*���rB
�&��#0���{@�Css��O�TVdP�	���18���+e�̝9\��>d'aZBPfa�F�ቧ���ۍ��g~Y���o�R��_o�EL��U~�
����13��J�I���`8��m��d�M2���4n�����?��3��᪭�cL��--�� �(��v��N�:Z/�]b��A}���T����x4,��1�u�˴��@3�6�~Ծ8Aϖ�T���
�N��L�2�Z+��%~ߌ#��aK��y�׸���@��V�w���V�L�b�c"q�$�-�n�&�m]d���,�A�w���3f��\�4�{�3����jɑߵ����C�K���3׬�rJi���Y4N	�:����p��&#��qlR�F��e'4^u�n6�^�>�E9�/ �*��	���>��'���t��qL�:����y�?=3�<Oҏ�d�̣���}~���N-Q:�r1��Ѐ�t�lE�݋n<�:-���EiY�.���ULm�w98��敶�9n]��4>z�4�or�t�<6UԊ�ʷ�і<h�J+��bz�w��y��^�2�~٬�#7�o�0�䌘����$ [���*#T��rRk�^?� ��៘.Т�eʼy��s�!�3�Q��B��D��oW��VN��]`{ٽ�rDXX�UP�@���:���-���p���A
M�ј\򞄄h�߾�2Qܩ��qK��\ �1�0������jʦ^Lu1�idEUp���X&�Zs�|�a���0��Y[ϱA�TNU���rx)x���e�Սq��Zshcu�{�:-
�I�H
⋉UX3˨�XV��Q2x�R����s����߇�ʗY���^_��D��N��r �N��O�Sn�Y��'U�~��urƮc��y�s��T_�nN��m����U'�\C܎c��}�0g����C��#_�������(��?"���������$����r>1S�u�	��V��W���#�`3�M�r��_�|Q��m�!
�����q���>���^ͶjiTާ�!�cS����a�q:z�!E����P0�㛇L-�X���I|{[#��&�gɗ*��@���ގ8�����
L�mv�z#���?�߮��*D�ا�T�"��S@*5��՝�҇M��;��"�#�-���ҷ��[OG��!��2sݯs��F.݄ p ��Kҋ3�pk��N�+c�E�p� �r�)�{���}����j�w���ŭ�0暑�}�_�[�w�+��]<e�Nƕ�	�6O����[��ǦnB�����+ۭ��
)#�P;K�wC9�=�s ���V,��\A�'��f��^J�s;��>!ŖA�Mx��q�\Pm�3�-P�|� $G<�3D;Ƿ����|/�T����a8����O��F�I��Z������I�ȶ馛Ѓ�v��(�͞<mj���~�2vb����Sb�+L�i'���n*5�!(�P�d��=��?�����ݸ[�9y@v�Ĉ"g������K�"�� X�[��ӟkb]�dv��(m�B ��NLr��U���&���V�l�$����@3t}��Uݻ4��A�VPQ:�� ��d���5�<���C� �Qn��H]�p�uY1�x��x������`�W��&�;ѼQ+a�Έ�AW��Nr�7�Lj�/�-tN2��֝[���`����z.<ӿ��z�}.��{���Qx�ym��W^y�OxQZu�c{P��g��o��6���V�M�},w�yq�܆�K�}M�\�5	�([�NȢG��oxyU��:�6��pɶ�b+ρ���/f6�o1U��r{z/�$��|�П��|����0y*�m�q�2#:~z��iqj��P����m#K���Hp���ɑ�Rլ�n�Sƕ: �����0�ZleT���,ְ�_#dÛj���lLi����;L�.䣮'\�5&D�M��$�I�oNƯZ��^{��*�4�������L�y)	�W��u���H��!�Z;�Wn���r�=O>0b~?^9��*WcvG�4H3Ր�	�qK��I�g�!JB�=|��y2��MU�C���W���1�(��/=j�N����C�N�/�yGEZWC�x�u�;+�Qnي�!C�찞�m&}g�9@H$�L�a�:���唼�����L ���qfՍ	Y ӳ��r����d���u���exI�xqK�z�N����S��,t��y+;��"h�d����	5��ӕn��f'3��4�A�G���?I�ma�+��=椹��M��7Wuq)��Y�PT��l���/���o���7�����k�ql����s'�W��bYk[^Sa��l��e"�1,~K�~ǒ�����ֆ?Zr"�p��]]���-^�8���-��Q��a��R���C�aߣ�^OO`ҍ4�){H)"�-5��Qu�sePY��X~3I���ϐ��(t�'��F��G#�����USK�0sD\�� .N	'R["�U�^7c܋��xI�-!���cfp{p�>I�edt����:�>MF�"�k��"���$'&S���UFv�fP ����5� ���B�Լ~���v���ʽ �C��1v�\����\/��w�����h��:�$���,M�2�,%�ϙ_ϛ�4�8#����G�E�Cp��-k�N�S#P~�&�Þw�l��@�x褪�땻�V6�c_��-�W������q�[ȣd��D�z�3y���[6���b V�6���G��W~�]�/���<��R�kwwұ����s�4q�(��{���O
��i��8�T@�ڰ�C5�^Q��q����D
a s|ܯ4�I`I�Uԫ��E�����N���I#3W�C�C�Ʀ�TSa?�o���ǁ�걁��:��[7��r�iY��r��1���Ѧq�.4��P�+z���n�s_޿�=䨾��T��#ҟ��H�X^M6�lg�:YMѨ�2|:��\~�c~�;*
��ވ��{�`������r�r&kN�a!��4�M�ڊ����&�T����xa�ȧ:SZ�#x�`�֭�Oa����>���V��K�_$7�p�m�$PJXG7܆�swJ�Ηx�'P�Hr�N5q������<<�x����O�sIE�*wжHfX��>Z�n���CP�����l�b�����ߥN���z.���+��Z�kaX��v�H���o�!�����9>u����z�ҁʫ��Y^&�3W��@0y=�&UY�D��q�2T����GZuxp{�\��� ��sH�1|w\݉��g��J4mG��n\��20ƙ$U2����D����Vn��Ƞ�މR�T9l��׃�M_�:Z=~�,z-�M�'��B��t"t�
�a����ۣ�^ ���S�5���^���ԲԞ�z�1���K9��P�ٱ��%�������*'��<��j�������$�t)�?=
)�.�i*~#nIyg�+f�d"�0�'b��os��7v�xo��v��v�r����H���c18w�U�@���@����O=>ݳ�?�=�����ry�Q�C#_{��� K�(���]	�r��t�Nr�) -��h �5�!�,�.�$>�P�H��O<�!y���d���#W��ՎJ�$��͠)��c��0��g�d��GH-=� %�0S�HOJ֢~�*o'q��V�?M���=(�%�g��k%4E���=�9���R@Si��o���I�`��\ U�ȸ��`O:�3�IfZF��Zp�F1��Զ�/���NF52'錋R-���43ڗ>�֜Tv��@2?��+
�F/��`�z���r���IzB:���UW�����Fg��n�"��f[����kQ�w�� ���}�a$o�0-��˦���*��B$6pE��9�a��~ ���`_�&�&�C�eS��:.E�tw6ݚ�M 1����S&���|CK�ޘ��/�N��"q��An�e�ǌ��ז�ǽ`k��L���B����=x	�8\��A.��B��RE��>i4
.K�q]�T��+Qm��E �z�1gx��ۿ��d���XS=��U I'��YZ�H�j<�:U�~ɽ���h��LTYU���m]��u�����_�D��3����C4|�wa5�3.�&e[-ʈ'8V�ɳ�Q��92
�e��9B!Ԧ3� oE3 aqTP'��G���1a��es�l�d��uA�rb[OC<�ٌOӏ� ���Űp��v��\0)�� ubX�����	iu��5�|$�tU�fqt1��,~�mH�	��b�	 ��&�ĸ�v2���5�y*$�������t]���p���3v+D+5D�@R�˪��C26G���l�#@�7��t�m|��,�N1����G���7�?�rQU��}�^Dnp�!z�3*%�w�˙5�����7>��=�J����#�2̡G-EsL�r���ogY�����@��/����4Sx�n���B�7R����Aj�(�L��g�(n8sq+1�dW���3:`��teedR�ndp�*��MD`Q���	]���y���5Bbv��l#��3Y�c�F�hx�{��C�K}����B����B��`/E6�pBS_D.k��zv":M� ��i+�+17�ֹu�C	Fi���"�5��t��I��Q�������Y��[�|�(|�Ǎ�`�v�;�e>�hS��.;p^��z�!Ek�л��������a�ɩz7�]4�5�'�rN���-��fW��(�i9C�!j��S�"w����A�S�R[��T6����%���7v|Tq�|�X�� Ϻlz�Ұ�y�h&��uԺvmK��W���EÄ����Q�6ޱ������Iq .�8A]��jw�ðTr��h�w�F���kJ:�鋻�~^A�'^E2�l�-�a��t�χ�xҔ�h׍>���):�g�Г��WY��#�,H�Oe����1�9�(<�yH��0��w<�6�,:i���-��}ﶾ�t�<��A���0<����I�[���T��?�>k�Ui_Dq%��>���W�}��v�.��AU�C֌����Za�=�+%�Qw8��srz�[o��� ���H���t^̻���wJ���t[��g]O�wV��DK�=��Gg7�;���/��{FzC��W�=`凈 g�`��1`
��W=�Kd���
K�ϭ+�t,�rD�(��Q�[s�~��6&S�/��
X&wwr!�W/�	Q��t�8������c����.�B�|vUt������F �@:>S`bř�qI.׏	��Pm��P*h:�0�J)��gR�����y?w�=s~����)�!\
銻�:����q[!��!�������@ʠ}?Q ��#2���կM��!�����I�	�y�������o aـx�Epc�g%�-�
5�}�K�JE�B�B��e}��3G��'�U��o�$�_oNZtM�{�~b��>����ڣ'�$ʢDl�Xx�_H�y�1e��FN�Q��Hh�mg��q���o��o�h E�.�Ӻ�~�*���_f�i|�}�$o3s?����h��0t�C�������b8&���Tҝ���k������"8�e��R��=��3	����=��)�{��HWQT�$��+>�&u�uE_�wz	i9�.��Kg�I*�be!���o�s}!�l�e��.�BD�����K��\c�q��Eiq
u���d �4��R��U����1�����g�� ��)R��K�����-��~�&f9����|�0��ۖZ:�}��t�;�51����S)I��D�p�jd�O���.[b9��HFOqp��־h���+�"y�����s�j6�`zy�������V�]~?���k)/��\?lԷ���%�FD���+OR#D:	J�hG
���SH�N����D/w�cj�p���>5�9���/�	��F�_51�_����n�-xE�mm�a��"?Pp�ʻ~5ͷ�~N����%��qFq�9��\%�-�@	h�R�= Ro��g�w�ZY^�����q4
_� g��ó�荁/Zl�����'���g��Ԑ�Y(�(�{�-���%Ek?*5�����3���O�[�v�>L��5�y����Ա��Rb��z�UЊ8;�1xs�G�5��2p	_Ʒ���;P�o��~9���;����{���x�苁~�w����Q��SR��k� =>���d�G'b6u�6ĲZ����׭r�>��ݞoy:q�'���댮�?��Ɩ��-O4��h���=ξ��\@Ԡ��}n�	U�:䨭z�E^�|�RD�Kd~m���ᩩ�h;�5�:T,�Dm��>��(��|ح���͍5��2vSbQ�j?m�z�8e�*���h��2Z�+r����	;�\{팺��׽�[N>������}z]�gO�~�̞�f75���.r�cB+���@4<G(��P��-V�×���ϕg<J��Ҹ�~�Hc�-�h�d�,}t�ݑcBC��A�B����K'b�L����K	B��Ӱ�(��� O3U���!�pɄ��cLGf{ ���b!�j9"�z�~S��L�*�	3���Sܥ�܁�j�rYQ�<uV0̀�/�Z�Z��Y���鞿z�@�*2�j�9Ͱ!�9�???,����#T`�t���sl��b�LK�̍��P<�`�(S���i^���K&e�k�[O$�Y5��T�-j�b����Xb��ʁB�KJ�.tC1yp�6~Q��R�$���8�bF�����;��'�cvqv�S���DY����S\�>��^���sD��s8�`���� Ĵ��GY*���(UV3������������Z��u��H�����p���4r�u����V�+�"�M��Tr�������Q���[��>\��d�@�¾��6�(����8wꯆ�NU��_�(Z�=0]cg��%��P�BO{L�|D�eN	r��Y�cx��&&H�]}��.o��?3���o�߻RD��$������]����n�x�>�C������!��)���(��13�����6���,U{w?1ݱ�:��u5Q�pi!},m5�!�J����)�Vh��"��اC�-E�]I�>��Vz��ܙ��Dɛ2��{�����~ �L���b����u�
� ��*9q1!_!y��������9�7�(��x
X^���	�Ҡ�i���]k��Lgi{���5Gb8��u���ܕ:��:]��/�����L���i�4�fV�,�R��ͩ�m->��o܂�+S����|S�6N������q�T�4��u�4p�-���yy��9���"���|��6	��'D�1�S�Y��|���$a�u���{3D[��[�'�>�<��ٝ��2�짘�!��V��~������m�T��E;�j��K��-�]��'��+�BU��������%hߎ `�f`&?����L����%l@�
�
����tu rQ��x򾼖wK�ȶ�[H�(�cn�JS0v���
�f|��A 쀏�SЦ��I5/Z:����N�_���!Kn���I�6P���\	���E�+a�dEJ.���u{��,���yR�u&� l�;g�qR��B�G���/�&GI���ޥ��B?"w�%b�;�<i��P�裴O���09���h�ŇLFM���(����D�S���RԴ<��^�b�c��*�Ui;CmQ�P�,��'�����(�{U�/M
��C<3���*�B�9D�41՘d����I6v{�bj_��̯��oL�,�Re�]�j6�g6�j�u�Z��op���<��N��\�{�&����.�p"�;n�߫�C,�h��%��	��o.���MS��,�P�Q���	_焸�.����i�*�!ֺ�,KH8sh�@�ݯp����0���Y��k�wX��P4�Wr��@FMy]23�1	9�v��� 3���#Z�oOs
���(���,=����PfF � ���5=�6Ӧ�Zi�)���+lؕ����1U��9��
��.�G� �4�R�&�������	"=ws{D,g�����8��.�p�a^�5���:�b��D��$[5�ǜ�zy�;:t�0����%���v�����7��Z�u@�q�]�'�� �!08�\�8�qJt�3���L0�Z|�%�c�a�w�[�(��VI(����
c�����݃�2��>�2Q�K�����U�h���B��F�֧}��m�R��a�V9��K��s)���׼{!{�X��&%䙳t����z?W�y��#��]��a��F�FWj�����U�T�<���u���P��k�n�T`�*�N�Y�PphF8U�������-���3o��aUOz�1�gU��T؋FY���p�k,����+��.@��,��s�B���]Źpz�2s������̻��6���ׂ,@�z5'[~��'W�)�.��7�WJF�hR`�RY��{���f�G7 ��tO�Cg�9�[����̭�l�� �����_�}�[��o�������;J�o�!%�����f����wwl��VL����X�0vg��$�
I1�k����7�2�_�P���U�1���70
Rw�{��`�矱:���@i�$K�.����{z���bdIe���4h�=~I�Lp:�H������|��T��G�~��t��h�@���B(`7� ��kY ������KMvL]4��7�x�3�b ��b�q���3��@��F�����>ʪr�b)�ݰq|z�p�:󏤝�WB���n![M�{r$ȾZ�Zі�z;c3�d��O����߶��S���N�9�?ObD���+�9���e/��&�$ð�]M�v�H�8�^�]#*(q��6=�R�*7w�ڟ�*��������䖏�Ҧ���4S���v>��+n��I3��]p6����-���^�Ϭ�T��0��y 0u�; ��9j�_7Zy]`[��)�O��0���\U���k���O1g\Б��%�HT����m��S�~��y�
��+������CM�0p
�^������Mr̟/��$�U�	>0�*i�q#�2��M̥g�0��s�h$5�K��Y&򌕯R��6��n���F��#͓K+W�?t�k��Ԍ����QY�X�ʾ���]}�m\bK���Y�nBD�pw�,�!:p��N����"V��0�J#�n��edX�S\7t�9.��r^����Q�6~�?@��R���9��+y�3��jiO #��dH��ؐ�I�M����BX�na~:�<�!��ƃLnWn���p>��u���J�b���#�5�̣������
��I<_�D����~DBw�4'�8Ķ*cГIը���~~��*�!k�N�`ЭhF��y-&'�&����S�rp�?tdZ������o
u�v��'d���0�0��\m�}�]�Y�W\��$���Mf�]��u��k��X��O���F�x8�uVa�����E�E�A�:��#�+��-����SFCa���� \������o|������ne<[Z�<%��!"���?��כ�Ym�e��;�� L�lSO��EA�����8^a�'?[��c�^C����:cMH����VΦ]a���n���j0aR��Y$2�
�ާE������y�ʼSd�j�-��z�@�q1���&�*�?"o��&X)��̴����}Tv�_���t����Ե3��ڣEJ�����)�'{���t�8gо
�d㝖S:�V �8셑K�~�0���"� P2��U_+�΅��e{���t"HT�p�F?Al���Չ0���a�b$q$�m
r�]O��Q0�`����7��b� ���釽*�:5*K�"���[3h�O�`�7	t�^1QXK�Đ�B{mO��W	ytM6�$�'J��s��MO	I���*�У����	 �YΥ�z�!���hw�1;,L0��G3�>ٛ/�I�Mĩ�6�둓��MEV��������3ZK�|�w�FKy9���!�rg+{IK�� �ψ+���}�,��6�Qf�)f��O�����
��xʔ��Y�$�:�{�@�b����I����{����k�G@H�a�R��dL�'���U�쎨K��P	��UV+{�t�����*J�8�8�����Ƴm$Jt�12�/��}r�|��T��c݄|QqWS;����\���	�ә��i�C�@��O�����'�?t�g�c��)-�K�ht�P��6�C��=JX	nBY7���Ŝ쵍��6�!|z�;EB��k�C�ù����6#S��-ڟ<��@��L"�����3��$�D�Ũ�7��f9;F ��"<7�o�؃j�PF��4; �	�2���	>܍K�g�3*<���?aM�Tab���T=��'w��.��G�p�{NM>>zi�-��c5Ru��{�-Fj��sV�/!֎Q�l��?`nϐ�ī+�\�u`���t�s�����̊;u密��+������87Q:*��5J�@O��=�-W��XǠP��x��c�q���wN;q��	#�a��C��9h�i�!԰I���^��%�gv�.�-�waQ��o���/��� �ܾ���<*;���Ψ@ t�������:�jE�`���H6����W��q��3Ĕ�������3�,�Y�ؔ9�,�b*{�9�GԏT��p���롬�\��MH��b������x��y�<2'�R�!ܯפ���`[�n�\��U� ����b��]	��z��g1D�T�+N-j���q}�O���d���)Z���읩$"���j�x3�M�#	d�o`�����$n�懮��nJ]�C��\f	����)��˔n�H�_l ���+�:	�v����8@��{O�
�q@>������[�u�Wԫ���f+CT�P�y���#���Pq��af����Ӱ�����۠�=�H��p� d��U�y���B����U=�""��ͺ�5�Af�[6uH#��h�����w��j���lr�0S�\������+�L�uɢ��p�q��v �w/��w�A�+v�&�1%��v]�H�����?Uꨬ9&���]�*[1ܘl��B�86��4����u��j�vک��A�[w�S����0�f.8<���BO**-�uSz@���u`?�~~!�Y��[n�N���uW���GWO�U�)t��B)��w�4���4�2�j��^�#��������8��\������a}��U�Q������:�e�)ȻV���J�2+t�V:��*u�ؼ`�B��yq��?W��:�V���j��}�|�0y߱��9Տ7�8���.<݊")J������v��u�`I��o��T!�uD(�ߺ��GA�M��/�Q�{>&���q�����jUf<����OT�%����̿��y��������0�.�K��~f]t}ą����*�ι�4��8�[_�D���
3��W(�ܴo[��J��&��(�a�;ƏDKj��/���#L�v��u<Ӡ�+���v���+��¥�2��i��NƤƘ�okl>*������j]������!��b)/T��l+="�.��(c}���D�O`r��۸��3�+�%����ᚓǽ��;�2����D�<��d~T��6��!'ͼ�6���DXT��V'4��W��ލ��[c2�E�HƤ�������/�{�w#�&)[>��܂�p�lIx�/g��:|�d�����CXw舻�3��Fa���>����۬��Ln�w���\NR�}m�)���dV%�+���ƃ��G�� ����
�k�
�%vG�h,��IR!�
.\6��j�?���3S{D�#���<�F�Q���7e�N]�U��"��
K���]	��a�YE�U!rLF�
�1�O9�)�eT���}����ת>��O������R�����,us�a0���E�P|�~5�eP
6)�)��X��.�zi�:�[��B\�.h�	V�,FƄ�r߯�y�;*��6aN+UCZ�P��Ҙ.�0���g3'ʼ�ae|�+�~�1�v����M]�L���hJ�s'y��̀t�;���n�	e���Qɡ5�Ϣ�cMW���<�+� �h�
dG܄ϼ�*�M�=J�}��Rֆ
((�E����Д��z��AήE|_�0Μ���z�/�34�/�]��V�l�X=_S:�ȵ�����fG��KL���)��(�O�7���2�5wk���L/|WGpu��2QH�r�K��Qh�Ϭ2�y�sR�,���rZ�,�f=�x�#RS|�W�gO�ȃ�������=�D��-�x�,�C�`o�#3�G�*_b蠀YpR��F��ߝ������?=%4~�Z�F\6�^;�˓��jL�Hl҃�O�d�43"b9���m���⼻XNdc�ַ�h�hR����|М�����ǛV���W.]}����Qn��8���od��t�X�'9��B%�|��C�s�>ہo`��u������TA�����x���t4�ݏeku}=��U�Fݥ�l2�:'�F󊂍e2����OH���/��C�Rm��l��,���~�]v���N�=���m��)���N�pm����׻���ur�q�T/?ԫ��8&���9�Dfm⫬�s�@�����`J��1�qǥY422��G ��.D5���J,!���s[����ٳ
����91�>�
1�?�@7��n���u�4�s��
C��cɞ�.T~�fe�����'aT����ޔͿ�����N���=4�t�7�~�n+;0ix�@���i"C�2�m�@�,:�[sDD�\�h
����sv8���'� ���#�Wz��Y���l�ېM�ᬺ8xe]�U�#�y�E��/ڎ"�7J���^�^�ً��L5h0�����9.�AO��U$p=�L�[1Y�X8JϬ�)���u_���U-�1�~r���>z@�������*\�0��E)Y%D�^w�Ԧ7�ڢ�: (;'�iHՄ����ܦ��47��I0]S������v��&�R�.�ۨ�
=hnv̓���b�$@�#�3^z�<���w\�� J1~PW��U��!�\����B��x5����ŀ@�<�X�� ��E7���}H�q�|������c��Qr,NY�����ٱB@[%c�ow����9���	�AO��/��Sn�͛q-	)�"����0i�[n���Q�%G?Ȁ1x2��o\���0o^Y�*������_OzK;��6th�@?Av��44ʩ�1���\jQN�б� �#o⯯�$w�"���.~5��:z�U�W���4�)v_���]���F�e����{�x��R��E����6��'���|�54O��M��D���ڞ�*dc���h��t�0�㒳:N��6�7!M�)F����^vu"f)҆2��$�L<�g�7(|Igi[ҁ��Z�M.܅k��|�L����z��k��t�.�.{-�a���y�_��.t����yȲ,��ţT��_K�3�ճ��-���R�Ć`�e��޹����a,�B�ܸ L�!�.S/r�.��y� -C�=8!3�l�^Z75G8vS�0��Uvѯ�����1�8�oUn�I��᳍�Y�s��IK���l}�$�� 5d5;-b�A~ǜ���s<�	�*�i�_l+d��mݥr_�E�'0xz�-.v�(��+�a@�j�j�.嘄��p����c��S#�ȇh�ƮF:\�2Vd6T"҅P�SB��FC5�OeDUS�p�1���$���T4��2�Mխ�-P�'��<v(ѱ�j�O8ݕE����B6�95TJ�G`�X�h��Nr��Q��eΑ�3�lV��`��B�D�Z?��7M��X#���z�ޔJ����"<bV�itD.���׽�T���vi���6l��Ăᘶ�B^gdcj|�w��B9��E��>	��0���\!�un�A�F^���7�ڧ�K��U����R� �v�
)
hZ�?���wS!~�7�|�k*�9:@`O�akk��"�	� ?o� �㙧r*Z:����B�������l�������x�;�[V��M�s3Z��J)q��C����m���o�+A+���{v�*!�:B�8�Gw�Xg#�jG3wbp��2���{���NWB$U�M���./�+������l�biua��|�Q��E���a�I3���m� ;�����3��7Jy�I��c��T�g��ފ����=���Y_�Xa#�%^��
����	k@�
|�8�Ʊ:���@�EV�52m��V$Jc:P���+��C��l�ZWH]�k+���қy��q��X�O`��܀rQ|�ojlȲ�@p���G7��%���}�sCz$Ο:�~�D�>�Q���7SP[h��u�,�-�Ao|�<w�+�W�0�|��|��)3��~lZ%����U�����U]��~l��ȋ���,��`���ډ�F��3N��#� t�oߜ�|�$�c�H��!Ң��Sr[Ou�k�g�`VK�JT9��F����煉iH��{Y�T�{��2=#۽E��P�������B�θp�쵗j??{
Y�n�*�Ԏ&�7�i����3���R"r��B�'����{���M�k�d'�����ەb��I���k�1Sݡ<�I��ۡ5G�R�OT�-5\j���.�E��vᲠ�e*�G�T??%|>�B���u�x���V���P��U�7�z����a��mby���vXoԦ�u����-�>�M���?C~:W(�R)6�7"�>�B����ۇ�K>��CY���թ|8>��0)ڻ�'M8�/��^�$�T���ѿ@	�{�;|����S�-��Yŵʷ7Z�C��6���^�<�,���~�-+<��#-��C�_�'�_OP;��?��%�A��J[*m�{�b�l%{����j��I�1�$�P�xkVA��M[���#�o����9�s�y*��t�vgMrTh2�Hbm�n��A%gN:��o�L�^٦�*D�`�( -�W�u����t0��B
��⪿�y��$����Ҳ�@[��l�)ק-�@(��ꮎ�7�q:������y�)e������T����6�r76H��Y�� ��$��1�U����Q[�AO����b�f�\S���Ϯ Q�����r��G�����&���rܒZ[�~"�Ř��6�B�Tφ���	���h�B�h�`�?�C�Z@�����N��D���p�����{~�՜qwvڕ,�A�R�X�ͼ#�
9|p�<7W'_ִ�� е�v��h����<�c`������d��$D�������J����� w;u�Q��/ߩDe�}������P6�+��6|~`�S��3P��	�-�W5���gZl�|�)�9��ݵ!2?�5�9j�%���	w��8�jl�ʆ��������:��T���|"!dLZz���X5��R�Jq)��j�ى毠�#Fn
A�tV��@���M皑���T�| �UT�5'���HG�I1�T��^�"I���$ZǠ5��������_	���A��WY�#�H	�д��>�:��c�3�lj�@u�-'���^!���F��m~�nX���@��࿑r��X�=1�8��� ���������6�{H�{��\���,DxF
�Q@���p��O'6⿀��2��%
�}"~�T�X��(2�X��Ϫ�x�T��늍p�;�1 S�@&�L�IJyTx����RoAz�<��EZ�I[B���.Ƹ�ǡ�My���M�<u (Jo���b.�zz��Q(��?7��ز25��Ṷȧ696$:��ҳ�kl���=*>3-c�~d��|l��^~��rJ� �S���(�O��rR�5���yg:�QJ>�g��〘�����0�]yoq�Aڑd��DstsK%ɨ�-~�������JG{�l�I��Cw����im��٩���|�lWA����V1��)y�ckl����4�U
���I����1��N!a�V�7��ή�İ�b�W}v&/2�m-Y����H>%h �e@��� o�mY���tJ'���p�����g��nIUi�U>6^]�q#ZN������ᲐlŤo��`w��72-�:m��De	�v�؀סĔ9#��\�{xϤ����L#���S�t�O0�G�2
��3�Ouz3 �Q����w2�S4J�܋VX"G��>Յ7^*���+�BY4*���\���v�%h�l���x�8���J�l�C4�.1r�,��coL3- �7o���3YLE���ߖ�����pf
�}��S��o����_m�SN��-���﫞�^��>Qa��R�27_$��	R�v�o�:��ٽ*��v:��iFS����_G!��$��X+�2ËH.3����j�W"���i.�i���4�\��*�7 �
������	���t{;�hy�Q��`�Hd�Ō_m�4Ḁ��%�ɜ���k�Ir�6|۔�l�c���s�/��#�A� �c?��(��p�ڻh�t�!�|/�ռ$����q�z$H��D�qV�G��ģ��x�o�����~A��G�J�_L���,����w���D�#J�	˯�� F�M��� i�_���h(��6m�F7��=����1�Y���������o{|�<GI�zX�4j�^�;_!�jF!�q�rԸjZ1��,HƥE2T{�ST�9�is�A��3]��,��$�Q�z��NY��i��a�a++�;@6�@��I��	��z[�XQ~p��{qgS�o�+$?vɏXS�6sK�?���
7m1�l_3����L�*���K�?4���x
���j�t~w�遲}7�+S�)���&π8u�f(��j$���>��8ߞ��y��.�S��D�{��ӱj���_1D��kב��(j��ԣ�`P���_�9��$�4��#	_J�d"�1�t��x�K���ۜIa��U~�n%���3�X�
*��K�,�wD1㈨68�e�6���gWZ�&;�����{5	T����d)f�q9�H�S5��2��wL�8��j�k�і�#����t�n9AǦ�VM�^� G]�W!fТ	��P$6�h��o����k�C���	��6�;z�ԕ�<��L�PG����T�/\�6��g�m·
D�����G�i°󬈂��N�	mhҴ*�"`����<s��]��z�_���B�+�Ѫc*2]AV�`�U��@�(zlrq�&��$��\m�M2��9A�Z�c	G�)����>TC�c�׈^�e�y��Ϲ�#һC���n�ض���ʘ.w�%@9.�0�����V'�GuÒPo�YSf"�9��D��6)�_nl"@n$�͒��	]R�(eJ�goڷb�����a�[x��M�?l�K�.��uB�-RBQbK'��yd��<�Z�u3n�1/���V/9z��lt쬚��T}X;֓�E;\Q.2l��Ѕ��
F�y��m�'�ޘ���>Q9'���:8��!�s�����b"��R���39ުv-�L�.6��o$)l�i�����~�V����M�ն%"9�BU{έ2�ǲ�����[1��a�7���Iϑ�g���Z��la]����D�ޟm��]V��G��
����� �nP����E��[�?_��H��5�]9������ڂq&l��ķ�����7_k�x$]83y���	��d1_��ꁰc5�/k.���+7��w���k<�]�,_�O�/ �.�	'm�b�8�M�����1W���u{��LNW�>�8]��`���0�t�wl��,e�
�� 1��;]y��8��x��>�1��p;s�|_��7������$Th]�o�ve��������]$h���v�'ge깝���<La;��Y��V-��Ʒ�����
��}w9-�-�:��`D���ً�-l�iN{:P�^���jȅ2t��6�uM�q���� @e!�{¹#��e����s��U��
e�.J�;��]t�$j�v��A,��&J h<�{I���Ig��k�@��Yt��ݢR$�q��Pl����{�w4�ה��E��ɸk3��_������mB��2�J\���14\��=^N;��C{��&OV�_�0��v�� ����3!�1���߈����B,-�R�p�+�ϭIaR�kt�����އ:$�x��-�m�
Š,sC�O Ȅ_����A^�Q��fp8�53�������BHws�2lh����iJ�bs�U�$8[��6l5\�zl� ��Ο&lmÂfJH�s�/H�\=nH�2^����I�E��o0�1����V��/��o�[~���P�S6�+�c�v�	χ�3lU��L_N�ٖ�LA0��sTO�5��^S_�%�6�=�g:���i1+�ߥ'?pG��.�Q�y G�20n��]>�x���|�a��g���Aν��:I�����h���ӱ�b�ϵ�Rc,��E��r���;����
,��v4��e�c'��"ˮ����O�[vR#U�yײ5]�����H�HQ�B���������%(uzI�я�<
����_��CX^aHJ~�t�>�W�;�"��B||��̘F������4x�Ze�	�L)�	��uh�,+Ru�ר'��6���n�t�$y��1��s���k/�\8�u�܎5��9��m7��%�먲U�Dz2)�<������ʇ:a_,#Ž5I���	3�5ˣ���!�x���#�5-[��&�����Xvw���)��Fo�î�P��F_M���T��r����𤖸�L��N�E�}#m��1�q��P�b�5B������q��㻈�[_�8�&�	��t
 ���_i�U�f;�U��:����YY6GNo�g)�5�ܓ�{����`��L�3)~7�oݻ�X����J������qjH#����M�	�uA�_S��l�$׹�ئ-n�<M�	�b��t��'�n'���0J: ���pM��߰/d��|Q˧f�x>�*p�����3F�3U�����G�A����[�͐�������4ڢ=�lݓ@�`��-8+*��p�PP� dp4�G,�o�d{+��%�azB�>����v\4D#����>��`����-������s�cd�r���g���cP��F�1�w��I}m���2�M�����s�TO�����죣P�#���`�&��N��}wv�� ���$Q潉�V��>���oB:��O��Z���}�s��~v�l��T/�DUc���r� �I�k;4y�H��ѷ�`
�u�����5�s�技�gQ��!H	�q��ȫ`�5�s��:���D@�I��(~}�y�Le���6�|��M���U0��F��p�D���@A�&{*w:�V�~*8H��edB�/��3�^��nG�NYC8�^}�U���x�D���K)s�ЭK���|W�k�-tV�A�ty:��팥��ט��a����047�0=��qR�U nO�0`�Io�͔�P���>�S�(���n�Z�9�$
]�aUޯ��r��_�y�#nhne[ :W0Fuo�e�*��S��[�#v�60]�0�%Ӱ�)QP�kѓ�F�VpZ��O����`��{%>sñ��j5\�u96Q�\S{P����-@E��5^"�"[S�z"��Т�4��I����ލ=���R
]��Q����n٧Ӱk�n�� ai�8	���ڌΤj	ȈO}�W�3�+��3�b�O-����Ep��`N��f�0�I�����2N��j�v8���3�ͅs����Am��5�^D�K=�i���N�@��`oxR�w]:@�Q)��:�n��d$�G�5����X��(A�i�Z�^HY��!�dؙD�lb΄'�=����o��POz���lB�1����?�U����$��Ϗ�?m��)'_�����@�˼�rh(�"��~�O���[���TS6χ�l>:miS�8���`t��3Y�����W*ڦ�Z���r�o؇s�U~��Չg��5�$���%}�U����@�I��D��<�e��2�"��iÏ`�v�M�X��D���7�|�bS�'u��X�����P!C3�/��l+H� �"lR:����9X ����������!z����AF�%M��C�mFCtf{��;���U�*�	�o]Z�)���mCn(ڤ�g���C&�%����+AXMf��դ ��%9G�ƃR��X@5��^`V)������?>G���?��r��ݦ�`z�e��+y�2�/���m���_ȫ�z��7����zг���5��"�&i�#�����`��V��%�Oi�"�-o��X���Ȍ��?�3�ATV��s�oy1>����]u��Aiv��Nl����n7��LeW}� 5_}�[豘 ^�"M�>�h���LR���-�FJ�>�k_��^��H����Ck�E��n!��<�U�[ێO]��kE֖�镉��˺�j?��<!�B{���rhr�a�6�u<�<˝,V��a\`����5�*0�� �����EN�͈���ɕ�[t�i?I��� ��.��3_�~�*E�Ʋ�Z�@���^�Tq�ɆË�~§�q���4�'ѕ	�r�[ `Ձ���Ķ��m�����h-�b5�Gs�L5�̾%Ԕ$���<�H���u��~u\��w��
5]B�"�- C��L���4;�&���(��@'\����;u<�K�����b��;���p,g�������\{W9=#"n�j���*[
vRC���62ł��ᑉC�L�����e�Z	X����9�����%�T��h`��M���4�l�=���هy���QA��?������ʅ�:�^��k�����m���.s��+�ބ���:�J�l��sUY���`������K$0x��Ek��/���@"���\l�6�,ܓ�+$*�H��ffuC�Wύ+�9^�e�!/���\A�ʽ]$Gq�H��1Qz%eQ���?����x)Y���s9�A�Yi��i&񑯐������>�h2]���դ�[��G44gR�� ����Q��d�`�0顅�H�5�V�쐽����
@��h�TC��L��[BH7o���~������s#9w��"�����2W�$���^V"ْԭ�p8cG��%���Ƣx���U����7䢶K6��Z����JF�B�Xv}�|R�j,�>2���d7C�X�⣻��֌.F��[K�����wZ��Gx��~i�]̃�D�t�ʓ����oKB70�TKK��{�@a�t+6>/p$G�¶��f�H�f�O8�fr
K
��R�����X�gR�{��W��RT�Rܳ��K#*�!i����Ãμ�ݼ�ߤ{�hz�1��<I�T��Xx���_�k�O�6:�]���U�tr�>�5a]�_���$�m�������f�N�U��I�ȃom��w�K5�XYd��^����0B�'���I�R$Dh�Y������׭{���x�`ʺP1_�l���%)F�rs���VS�%���=�ZP?^��Z^�fǩa�$	��)W�k�GHMd��6ZY�%(�R�}<�ܥ9�3�.o�P����[+� %�B!�͋ .����:GQkc}A�A��1�c
Tb��AM���������h�i3���-O������Mv_�/	.�
���0�]�p�ؒ�M}|~V�|~.T��s@Q�������:8G�Q�������%���'�K��C;�h��v8�G���!�z��=tD�5��ϙiY�8qO��]��uaq�x�_F��$�e��7�d��鵓~�+P��<鄓�r�sip�.�"�-��({�u^e���X�:�:��h~��&ߟ/u�/�@L�6�sG�(�6���J?��(z�چǾ a��dZ��S�+��&�3�:Nk˗��P���~@�V�m��D����K�"���.�2��_l:���x�&���:��W�3�\%��Z��I�*�?��"#���PؤC��e�V5J���ĩ΁N�nge���ӹ���^'{�S�LL���N�T������9L٘����#�:ʜu*�q�cth ��`�n<蛂E��)Y�������2o\ߺ��7l���Ǜ����|��?f#��
/����0t����d�Ǵ�����7_�1�9�jªBP��qLӁ��4����i��0�$��B�~t�X��p@����]������$�0���R������/tg��q�K�	�3�T���?�� �����*�v�K���%����
?/ #_}<��
2�:~#�� D.���'�j��H"j���I\�����$$�c�id��K��j���]�%C}�]�IMI�mͶ���%���}ܙ�'������h�~��.��n�aѾ�e9�nKN����Q��L��3��R�D�SI��́`RUh�4L���L��E�sWA.}a/	�rc��"SB�E��x�A���`wP�h�(rF�W����']4H'�Ji-Ѩ^���*=��/<���-�{�9�=0,b��3���--���6��h	!.���Ȳ�R^<�?�6ɐ�H�m!ЯT�+'�ظY����UDxٵ0�ٙo#�9�l�U�)����o�B�K�"Fzt��A}X�|�K�y�]�L|j��@1�s��]��2�j
��t�P�el>4(VJS�a)N/./xv�}3Dc��A�&��48�U�V�׉�Ӻ����WC$�����Ų�O]/�nQ���.�3w���:���0��C�( ێ��� �C;�����E�����.�yx�>��8��U�ζW��g,d=��j���.������q3b��:Fl,�EYP'a��hf!�cx�9��J����iT5	˽��=))ʖn?�Ȗ��;����i����4@c��y�����	���0���،�)�����YaMtH{[�{��8*&�W���|S��|��]�eȰ��p^��4��YG������-C��fq�
��]�2"13N��6ȩmyl�7'_�Q��xi*-������na�q��$"�@��u��r�+��ef��s�;v�.�	ê !�*b�(nl��*�6ɼ��)&V���9G::$���9��q�U�_%&�v�E$!@�sTXL�OD��W��%�X_�]��q�����	ka��HM�E���b����пM&�U����ʌ?}4�6��]�
gJ�+�s0o�����o[�UӶ��xCpXq�s�IX9�$�a�5�@��t:�I�h�����ŏ�+��fĘ��&����ss�uηE��^���RM�����V����^J��0�݃rA|�����Ɇj"�J��_�[���cSpǴ���!]��^4�\�[���y�c4aal�/��^|;<X#h,��0&�'_�PP�Ҙ�'�r���pM����'܎�V�)�͟2QS� �U�Y�ȑo5T�\ /�^�Ҥ��@HSq��H繶X6)ƚJ�s?����ɞ�f�+��)���*�+B�b0�v���d�_u���	��W� ���<!�I�k�
V+�9�ek�� f�1�\��"%H��/˘�]�i|��R��M�"�/�jB&d�sS�Ca��� _C�6���+����;0S^p6-���'*��ׅu���Z�dι�� {=�#�R����2���]K���ypF��Ju ɋ�ߎ�A?�ud�� x+[�NF���D��n/�jU~Bb�0��0�65�e�l!��أ=���@YE㩮���u����_��3�/#g4:���y[��R��a��3*g��$}ל�y�K��+K��kn��M�p鳗%��^����i�jt$��8�i3�bʮ'�C��ޓ�#���]��Z6!>�g�\d�c27�Ҷ9�
h'߹ 8�[��aF��M�?<T�(�D2�b�kN3�M�'��"�,t2��n~ ��T����S�Ae
�8��$�ڍW�4�G��)@֮@���Ҁ�vu�Ȏ���63no�W�@57ǘ�WQ��s�V�X�����&��3���>�5C���_�9�կd�]MA)~�m.1O���b��t�O��"����|�i(ޟ������s;1���G�a���dX`mQhz3����uo���AI��=<g��,�S��I�N[k|9�^wA}c`������!oE��a�Z0b�W+��������<���e"�-�^6:V[)gV]Tm&��&[r�<�"��~��r�:���<z��?�n[����֋�V-po�lbY�k =�꺾w��UR��F���EU�ԋf�����f��ر�Q
��ig��>�~{<,8���O���V�&�<A��KU�T�à�_k���-�v�\��^�4�?x�낮r9��? �_�-�.�`i���aۉ8�%�*�o�I~%F��i;��aJ���Z̝��(�^��ȭ�����c��#w�)��SġҚ����-Uzׯ����r�n��t����΃K� �8�~����R=M�4��H���
2�c� #o#f���fB��A�fP��,�?VU�L�a
�R��V�w��u|��90�$�j;�?�(����}�x.Y��t#����	��'Z?v�$Mv q!rg��+Ch�Q� ����,<[�_�W��JЗ5q~!�yX�`ڏ�,"ɤ}(�#��L�W����Q��C8�.���&^��,�P	e��@!!��m��:�,~	���b���W*�f��E5ꔟ�Jv�����Y�M���J�{�����{8����%�u�c����� `�ye���A�e"4����^�%�K�����4[�~V�-���Y�zZ�b�3�d`!�e͒)���� �CL���tZ����obu�.}�Psa���g�C.��.���l�-2�~�
���^��K��;[��DE)�Y�۝#�Vׯ)A�#;���4r���1�;�ǹ�7T��&����>Z34��ۑ���|�pΰ.�`��o>�"cn/��F������蜮�toH����8�X&��H"����3��H���'���Yp�'�2��7�n�n�@�*�pxd�yE�j�)1gC�b�Sg]W��{긓�̧���c�)B��8��f:c�e��'Ɩ�4\1���V��T�JvBYMp������_Q��m쮷����B�����h�j� �J���Ä��Fa�c9D�g����zX�4�$̈́�P�.sr t4!��ՒN����1�kF�cw7([Oo�'{I���f\����s�N;�K��r�	]�>Ӂ�>TM�����O�O�d�Н]�5"�E��0\e����%˯wR����	�泆��b�Ҥ��P��ٚ��C��[�+�6`�0���2s"��E
v�6�>���=�G�.��@���=#/.�n[�H�<��sY�,�T��*>�w�(.WfD�5S�O5f��0��+�*-5��;�u��W�D�fIx���K+c`!���>@�;Xa؀K	�A��iW��"���X������2�X�X�9��v�������89�^�-\��h���$k���?��J��~ɶ8�BE�v��&�����v5"��U5�I��*��իjǨ R˷ �v'%µ��B^*���3m<*�tR����)�/�>��r^TP��V��{�V��v!�ռgh��3���X�2��*�����s�ę�
aT�f��^/${9m���8�~Xv:֋>`B:O��*��������{)(��u9���=�5����`���d�;d��h�������l1��f΁x���e
dw��$�0mk�ߓ�a�_�7h�����'�ܟ�6����}ͱ�-s`�jƊ�8UT����H��l
���S��O�5�O��r>��W1��>��un� �!A���+�j ]�&�~�F=��N��Vh!�۳�[�Nß�X�P�����C�~�f8+2�&PEҐX҂�K�[~���y�v����.��K9����4Z�\���Ś3ˈ�2:"�v�z@A��o�������@ǡ�j�������M���g�ZQ*MG�R(3�V�D��އuƼX��*�r�a�M+l�����yBђqI��#q��䪑&�4���
X&(���\AV��N�Y{�/�֒�`��&�gX�}~�E�+�]664�ڈk!�'}�*F�!{*��;%39ph�Asl��F-����W1eZ���)"#�ռ8�qkQ6ه��	Y�'�,:ͻ6����J���`��.;�ʏA���=R"���N���	f����/�q�qH��c�����e*=�;o�t�/��8�崌�R}�g �A_�Hy�s�Ӫ���)���%��A�\�o��2�s4z�b*����vt����W���&d��Εpw��UC�tO v�qJ5��D/�?kΤ����VL�&��͞��薊�wj5��ke'�Vd:zZ$�h=�h,Mq�.����p��N?�rz��*��N���A!����Sާ���ؑ�.w�l��U�������T+z	��7�x��K����+�Ҽ	2��1��i>��Ln�=@�E��7)�u��̕J'끙�2�ȶY��+���Y �vm���уne��i��Ҭ���30l�v�.�M.�rD`��GN���;����B���E]��f�hL�)�{n�_db�Pˇ~*�������n��Q{���9ScQR�i��,!{C:H�	K�����ք�-F�^ൗuLzb��2(&t��X,�� 
LOb]�\>A2~��`�z��̧8�|�v�ȃ/<YNb&�����u8����,q\e@�0'+�쳤�x]�m�E;v�����޶S��}�7�̢�_�L��E���۾����n�$:
s�B�L.�
��\�<}�_��Ib�$�ˀ���ަ�Q��>`��e6���D�3j���ꐷ�� ч���1��$���\@\b�P�Q�^���q.s�e�qD����O+h�H.���S�6�G�&�2�n#�<*��V;T��^v��o�,� 5��\�y��$�z05,�v��X�v[�PHq���S��ys�N��:����(p���Q�W����6���r?2��¸ϊz��ַ��lÇaU�&�Q\܏P9�N�����G�iq��=c�$ �]���x��)ݗC��R�zi�.��*w��r�}��b�A����΍��+"9��X����[��-�o8�2��H�
p��?�\��(���Ƀ�7%�u;��*>�ʤ��B�L�V���qlȢ(xy��dx� .��쌳��c��a�/��a:��iz�!�΃\oT ��w2s4�T��^uqm��_~�Ѭ�5��P��6���v��q6�w��4��-6UL�B. ʒ;rP��czW�R���^Q�p'_��F9�^z��lh��N��S|��l�ݙL@©�I��!�e�	��Q�oY2�F�1bf��:a�̴&�T1ý�o�oiGޑ蛢'%�R9�xM#h��P�cH,�&k�'Ğ̰��vw�r��cy��6�1�'~��� rw��NkKK��$�EL�''�	�q�l�8c��=���$��$|Q���\�{��n�����?h�����"���h�����r�,}�W(����Z�&"r��RbIe���(��<�n�[kV�:��{���j��T]�tD�5���fx�(�:R!]��!�}�h��/�-��uN۰L>8_�������U�(��Xc^evUS���d����'C�'#B�J�W^딛RlK��=[t_��Q��,�E+�F����d��+�g���L-��J4_G��F��1�+���΄󁭋Q	�`tv$��j�~��d�^�ifR������U	Ѹ�$�g3�_aEaɚ�ȝ�ƀ�"n�C���ԽT�S3N����0��| kU��.���V͒���9ܮ�p�P���br�����j�����O��t*�o���M��T@�  o�g��'k�W�4�)j�UR���B?����zK�N�y����'��"u�uB/ڈ�z�*Ue7^��P>�]q�]&'Y�p^7�z���S��Lw_2H��ZRA�|'Lb�k�y�f�5���{�v@��7������݉9�z+�;B�J?=�(�<�k����p��%�9�o<������$9��D$^Y@Q\��&`Z8��-��au�Zj�?t��E��te~�j'�9@�dO��֪�G�#ǩ..8�:��u��L��/�>Z?{إ�Q8��b~�ٶ�����ԝ��k��p[��d���+�Q�bXm�(�Y��\�5�ܒǃ�/(���m;��,	-�dz	Yj�뉔IȽ���߬��,���� ��ޞ?JHQqQ/��'��v�S�m��E'w�~��mc⌛f_ve61�׹O������R��C��D`�j>	�=�O@@�ep�EgK��]�(����~d^��q����.�� {�r���@��'��f��/{�2/�'��ڪ�Jbp���@�t��0� %�BG�K2M����;{�r�$5e͊@I��<��!�x�8������q��[mˮG�!_�th�g7%$��⮣
�u�n�{v2,�����tN��_Fw����_��X�-�MC3�T֍D��P�O������LR����M:�M���(l3�hn��b�}�S�kGȑ`j���G������Vnd!�SB �+��7���V)Wk�U�&�i�#�ԉlv�-�K�L�3��)1�mw}�ʟ�����z�|�تc0�w�)�Ԅ�C�����蜿J[̩-N��޼/��c�ջ>-���Qo_�Ό'kaV��U4!�or-�ޗ�(tT �L�������-c*z�����_�lX��qlβ��ff�<!�D�P?�![�I5�~-�u���;�D���<^�������(�������=HQQb������<����޺A!�ݮ�Ch�1�ZBsC)t^���93�p�x6>=�Y��+���K�m�1w"����l����?:���t���)�����Z�%t�
h`���'�-��kY�0�v��J�8�]W�U�.��7}�b�>nK\Rn�����.�]�����֖����|�s�Cs�4��-�l�<���Yyp�B
��lC,$��W?���X*����k�������y�8�Fbuٗyb��s��� �yj!�~XT��e�rj��=�`%%
����V+��h8�j�h����L�*C�	�z��&�$�!��{�'�.��f�e5R┼G�Z�J-�x���N�t�B�'���Tf�U�x�q_�ѝ�C�/�~�#ίx��oZ�����W�	\�J�(� ���i��� \z��},~W�S3D���_j�rc�ť�9�ר%QΆ�� �b�
/[�K�9�R�zu���ZqV����OX
�j��kwU�ťݙ�w\�3�����o��_�Xr0$�ȧ�wZ�V��1��o��o<>R~Ƽ���&w!$����-R�{ͨ���q�OH��9�K0!ز�s���IWe�a�c|�f�{eC���څ��[\sԋ�n�G�@�A�s��i|�'��x���s�o�d��y�s�aY@�Χ�*�Ku��yD�&@e���j}�ԗ(rO�s�` A�l�]��}���y��/:���7¹S�J;���$$��pn)՚�#�JE���s¼l��cb`~]�W;��=;�u=�7��˕��Us�ZVS�'1�iA!h�z���B��L�4p�C��"�EF���(U�,�1?�j4Y�ҝ��פKs.�М$���������e�s{���h����d� ����e�p�3~��?�[Ћ���	GM6oN c��������FC��M���)�geeC�����:�ѷ�S��b9�<��@�;&�����6�Aw�x��2�&�`Gr�\�	��b���b+U(S���R�_e_�@�����0��'�n`��Lq�Q��9��OIf��!�K��n���1]��z��Ε��Z�������%�T������ئ���`[b�(�`[e��:eh9���el�d*��*� F�EH��9d&��ms����65|��#vAn	ptK�p^0,�!���]Kw,���٫��ô�5\�V����1�7(=&��pb]�G'�b��OƟ����;����U��f��Z�I	��_B�W�����ԁ��a����I�SkZ�I��R�f�oϞh	�K��C�}�0��y�L�E�^�����䍝��.ig#K�r�	��kF8�Y7�	�t;D�튮�����d�x0zG���9�����	�C�v�б�qb���u5f$8�α/G(��CIl��T���zI6�o{�4��N)�a�>�g ���*�=ͅ��=x�>X���Ki:���؉iG�H�E����|n�����^bEZ�%l0��*-�w��Oٺ.��Q�[n��(�c�jcs��ܬ�T�n����&�Ϳ��G��R�
"!)��	FD"�Y��ҥ[�;�$h���7����
����m�w*`}�d����S�bLB�	�Dx����C���~�����%�SR.�>��9�g�}T�8�HQ��� ��)�e�=��tf\��~�6��
�&�Ό,�$���+
l;E���P�"�V����^1��{���s��F	�j跗�UC��(�����]I{�UQ-$q��`�j^/�d�۬�p�U*"��kB���Z�':f��,\(��J	�?��D�k#��BoJ#L<aֿγ��1�p��J������Z�9i�f]u��)k<q#%�>�=o6\���h�t���ۉ������'�o�@�ғX6Qi��i�6��s���M�D^��=�� 
����Ȍ1<˻S�9ٱ�����_�߮����{��:�9�^����s��?�xЩ���jq�̝�&���:�u!r���gK�5��G���aD�M��:��/[��]�/�1�<�$��z�4~F6,��Ή�i�)�Rφ�-C�_�â�tkF7��c7e Yg;�O=}���,b|���r�Qf�u�ՙ(� �ƹ�9w'��S�_�)[X�@ȃ�͟�l��ǥE��oȏ��d���40s�<-ӐP;�}z�d���3.B��@�F�Ml������yf��:h�@k*{<b��6�Y��풒��m�{?�)��Ώ�qӧz����Y�Js�&@�"ƶtM�ĸƳ��@�U���@�>�N��/ê�غb�Z�X1Fd���mn�a��_�HŊ�_�^�*a˵r�u�Cf��h|@7��Z"ZL-����b�M���8�"أ�pX�<��̐W��t�P*E !8���F,�'Y�vAr������7�h�|!#��v��o$W����K��r�?
懹�������i>�Ⱥ�v7�.@�@��8���:
<EQ���D�4�!d^�~={I��(p��n���=�F5�6�K� ��F�qv��i�22���bO��S�v���g�u��:Z}����B�����X}���z`_�ľ�^��c�H��d�5�M�j�&;�$ę== E/��y���6�J	g� �#��E:'�c�<S�o��@��Q���o0ym��˸W�Ĩs-�%0��h��Y(���ԸvS���.D(��H�#��}$�S�Qt{�NF}F:�I�a�y|E�����QN=z�|g>zw�A氘\�����I�a��g;������f��ޤ�4P6��d���ge����~s��V���j�ə�̰�t?�*�f�災yX��&|s�Ų���S�L6_y��]u�������ݩ[q�u\�z���N��S;t�(8f���s�Mf�����2�l������U���Yb���у\���~7Y���KU�D�d�~7	(*���d��K�g�-nK?�#P-1�-��lj��Vk�OR�������q�[��OpM��u��+�ab6�x���gN�,���W�!��
J���+	°C���i�6�R��-����銚@�����T��۪��)����-FR}ρ��X��L��.��(��R��/[")#�3}�[鷖��9��!�O���ǁ`*�aKz{(��i3��6�i��K~�XC�@͟����+�F������C������O҉`V)vxA���u������B
�w'i��a{�9+Y���>-��M6>�ěv$.�`�;�K���j
q�D�x�tHg���s ��� ���Km�x1}e��]���7�эI��c	-�np��jU:�����4�G�	Q������h'+p�v�%�2�:���y���' ����������nŝO?����"�CeC��z��+���t��3c�C���Y�~�J(�Na�������t���HO��S1�Q�8˥��!�<]S�vP��·���=Z ����C�;A�씖.DV��Vٟ7)i�����s����7������F�	&&
(�|i�j�]�4N��3Y�c�԰�"ޥ��3���K���@�/{3nΉ������#�w� ���Q̟���#��2u��w�~
�AI����{�Ɓ�C�R��x��؂�y3ӥ��чѨ"������sb���Y�9���TxY�
��:a-���^��H�����u��(��	�O�j���Gc�1:6n��'Y\��`����B@�n�ͥ�F-��������Nhξ+�bwK6�N�-�F��@-PB�B9|���+:��%��7�q#ޫ����5)�O�t��7�M�N�lŠ�1Eeu�������YLj� $]p�g`ݒ��[��H�0f1"��Q ^�2h�3�5�P�O^�6ao�L-�YU����9M��m�f ��һl$) ��+U`jvp,P��D�r���$� :�p���Ț���n�Nީ2�Ȋ��i9:T�z.�b���>! �������!G�v��ڃχ�"�)̳X�E����+�:@s$֔��\�ጐ0/ui�'��iȎ�
���h�Ud�dcAڶF>#c�q�43�����f��2�*b�q����tC�*p~��{x���y��N�!���?M+A���J�����>ZK>]����~1�g�����ҷx�z��i`��g�hٳ���z������/���WΘ��Rn���(����rci���1��:�M��	��E��WKR��*`������}�U��W3�����;������s�K�r��l o`U�[�EE,��2�>\�Yز�;��W=}X�����΃C��I�^3�4�T�
 r��{���c����C'Ĥ�=�͞=4ϯsƺr����͈�t�/©�4��.P�I9����4�R�e�Rx��z��Ng-��:����Ȝ������tE�)�F��_t0WY�} 쯔�LL{v%g�$��]��1�n9q�|��	h�_2��k�F�7��c���c2�o��|UB(��9r=�ޥH��(V��]3}��G?V�\�dg�c�[���v�,(=C���I�N�@�J�{-h]����^����I=����?��2`�j�Ar���+W,�Xr����xPChhhX��Y��<o�D��E����4?�k��Y�YU��ZɝrS�qJ�$Z�*�`�:wI/�h�D��Vo��d����P&�d5�5$c���6t-����ȶ��u�؞	_�`¡/@���gߏUr5��Kyܱ�~�%��g���48F���R ��蔕���Ú�=�����o�Iި�'��@�	��G�#��l`��en��ݼh'*� �D����و��_���P9�C�U輭�߲�I��Z��O��0����h�M"S�e��/��^32���9<0��L�U1	�0i��,�su^�f��|5�4�J�������5�vgS�L>Y�~+������!�xHG���7o�0` �xZ>A����Z��'�jյY�@��Z�k!JJ=�X��X�Ǎ���y/)0������콖�E�)�f����
k6>y�b.JuWԈW��M����<�9N�&�T\�_��$�9>��9�oɟ�Cc-K���$�ԄI���	��F�7�- )�L�*���!?5�-�����\P�¼f�_��+���kA	������T�[�kVǅ�7�8D9����)�{X���"�d��S���t��?�3�Z���8c��XEe�]��)�i-ʿ�*��8-�]��_���a����n�e�s8w������A"%ÖM��#��b���l�H|�Ǐ�g:Z(5؂�I�>Y^#��?h=�8�5R|/T�ґ�-,y��|#��I�jE�4|:�~��y]5�>RQ�H�:.��1F��=���x b��w�촍%C���YD��-�[�5��y�L8;{�ф���w���Ȣ`cVs��|9ӈz�yyX�,��8��k4v�D6�8^<x"�q�b�L0"��Ծ�>���� Y�PCR���6������r��}}G�������1��3� -��
3$[�?���Y��Z(֙ �n7*&l%��|�B�1��9��	���?R�]������+�hX���^�N!��¦���y9#�	o�TN��5Q�O�������0��9�X�����O�%�p7�'�C  �YtA��Q�ӧe]:�U`����7���M�)�Բ%��2�i�Qo���!ԣ��v�n��[F�q�H������>�NR�V������7/�阛߲�Z�����.Nax�@��Y��5��֓��;c� ��,f��ў��e����� > (63�X��a?���L�N��5�g�@x��r�9�w5�ݲt��q�5�����3���m��8	  _��/W��M0�������U/�[�)�߸���y~�Pr��U�-&o2Ʒ�u\����J����!F{2RY�B3]� ��AR8s�v����gV���t��Xl�!�RFQ��%V���cr��0+�����B����?!�~+�R�����cP�?9o��;�J "������^���T�ua�[�� �RMp��'D�T%X�{5�|	�z��r�G�?r�p�W���ٔp$�Ϛ��� ؄��9��/a+�^X������D��.����Ъ�XGWU��D� ��x��(�źM>],�BP-�|x ���.�8�i�9F`?:]��h����#,EY�i�e/Qk��)r�17㇦.��k��m�:r2�~�A���¡�A���7�o�f��պ�F�����J�C`9œZ�\U���m;H��"���I�2���@ܒ��k�`�l�L�J���I�
��'��Ln�9/^��37��;��P���6	��/�I��uY�U{.�.J#fm��G�mwm��ǐ��o֑El�u|���F�������v�{,>[U>�x�~N�� ��-�g�!H����mn�55�ysu}4��!7|H���<�v���7���)�-{?IbPq��Z�{c��X�ռ�UQSO�(�`�&�b�u�TJE���@?���58�$1��I�X
�+��O�O D�bRHH�����\�(@���[��V��T0�h��ȈI���^,u?q��cYu�;>ax��V�*$���@_�)��:蛫���2���1�E���{Ff�����������M���!���+* ��3n��������fri������Z��6�jw�`����PAm�����ʋ�=ߓ�*^�K4]\�LG�\/�jb�wn��#�?;�K@F;}TP������t$�|ݚ��+�OQA�����ҋ�ٰl����H9��2�|0=��(݀ʯiu�&����l_�ݲ@��(Yu��B��r��@�p�^�d޷��}>��yO@4����h^K4G��4���_���[#Ǣox����*w�EB7ӯ�~f�c$�+I:=�|��o|���̲��<��^2�3����fi������8��������'��VQоU�Zm�%B�5	�X��U�,{?+}��>��6��6Q�����42���;�����.�;"��V"�ڴ�)���c�4�7VQ
9wZ&���.M����=$2:8C� � ��]v��k�7N��m����i�d|Ӡ|��ش����M� ~j�55$�O��H �w��*��צ��h�&��l���*g?����KZd���q����%��z�+����디����"����ȵM� �a:��&��x���HAS*�`�[�V��CU�$�
{{o�h:Y����r�
���u_;#�HNۧ�=A�P ��5I=�S������5H�����eEgZ� gK�d@
Xce��\$�| ����-��k�Oav�1'� �֦��~l��-�'q��;��q�o���{�;S�i��t�˥�5�o($�ҿ��Q������;߷�g׈,IC���˿�O0��2(O=
����Du3y����,r���=�p0�4崆6�0V._��j8�vox���H�I��C$ʅ%��ѣb�`_7�͢�}[����{ef�gy�
W��-&�8���z���ʳ��o�+m��ε��G&�(������^
i�yR�;��5�;�Z�$%3��?�5%F+"�?���t.���q1E�����&�^^.�(�����v<E��8_�F�b�W�hK	�&��'�b_o&������7����J�AG�?�m��S�@�= \�k !�2�T��&#��B?��t��:��@z(��\��ny]?�Y��D�=�pc[���<�KZ����u�`/P��������\g��-����uA /���,�\���2��p�!�Ҿq-.��a��vʺ�����dǜ�qG�b�S=+�-�}��0<���7�+�H��+�7YQD���c��G{�5gfK%ہ��v��X�?��lď�1�����QP�F�1�M�Ӷ�7�?�A5pw$L���4��lD#�� X��O~��̻W�c���E
ɷ��lx^�����"j��H���ݨ�U�����5>��h��>�]p��f�ϿS_Z[���*]}�#��P���$�
�����;[�ĝ���g�]9乕��_J����;�X�ܗt%��M�b/C2v#j�4M��`���B�2��(�澉\#]�� ��#.�wgz����QP8�W3q���VGݶ����~WN'Ox�۰I��l,?��t����P{����}X<�d-�V��HI���o-3�~�#��\;	T��e) ,�.�s�G�ڦ�L�E�u &��@��^a H\���rFBmZ����@�?�I Mw�4��^���p���pK�����ug��ִ�Zށ� ���T��|�����˺:��W�4=�4��8��*��A�J��I�L��a��[y��-d�����4�$��t`Iݚ�Ө�[[I��!�r�VH�X���ivy��h������Xİ��"�D��=�$k��]&^�1�>Rd��ⶸ���RzkuTZ|���$��M� ��	>����y |�"{�r?���W�9p}Į���*�
��Mj�*��x��u��`ac��/����_b$'�U#� ��&<�%u�>��s7���Jn(��(g�>�0�Gr}��d5�n��k��⺝[%.Ww���n?�˰;c:�Z��u��T?�c�QC���PȺﹳd]��\���,G�yXk �4���� �F�L�CK�x�N�q`+h3߳+��ֹ���x�h�U�{�,7�e��腘����zT�.\���� u�����J��1e��N�0`$�|����Y䮂�4�v��Њ�w ����&5�����0v�pS�pʴ�G�n��`v�����t~�#�&	�;��<Q����f `��u�"�ib��f���צ� ��|ɗ�A��c�����#��w��w�;��[�tk�cV�1��i^���q �[ݭ��6۸�������
Onɂx��X�vA��LHDbs�=tq͵�7�p��]��-JY��[���u�D��5��`"��wE�Ӟ:�s-�ߥ��f���@g�a#��`������_9B����Q,/�-,�����?`8��u�5p���ӵ"����LG%�9���u�(����F�}������)���<� ��_A5-UՅ�X��gD���/�5�Zm�mK��c����Y6��~@<M�ޝm�#P�L����
��IE��o�?[�o�x�<9#�tMfr��"L8m�te��� �&x�)%�g�@��$B���4�sg�$��>���6COJ�r,F�Z)�ſ�~ �W�)���g#�.��F�t%��h�#�������G�vQ�V��J֧�C߅6<ڿR�i��vSE7["��p������d�D��R^#/�辨�fUf�m�	�,@�Ы+k��!3i������N�i���>�hp�c�i^qcyo�ľ2�B���Xy�!{��*WJr��(��tYx�c-s�Ȅ|�η܇��|�BN�\~ �B����^�x1ae9�qTrc��� ���<L�-��VZ���ES��J�NX��# g�;���w*�v+Q���=+��iI�m�p��sU�����:��$�~�e��EG[Ux��S+��E�7�9�v��;��6�3�.�\��;4.��J�Q�f^���KH��Z9fT0e�jl���[@f�����9�k;�e�H;a�j�)(ZQ�H���dd�vTi�9��#�K�dE8&��͋�����a�?N�_'(�NC�����n/�䤌e97͸s�&����F�H<����	��v��!�w��L��o�y����~(�����u�t�V����.���'=����E�� 5/����`lêD͊Cz��~�{��8� �psT��ſ0�Y�Dp�v> ����<�'�\�p=�~�Ѷ��iE�G��U?(ΚuT�=�Zn}h�	����'�M�����A夋u4w��g<���{��2�߻�q�b�:��u��h���ڨY�yH��+fb��!����-Ut��:e�k��'������K��ށVQZ�����!���稭�)���d_��{�/������^��
!˅�u�I(���������JS,̹��7NU�FkN��]@���e.Q�����%I���*�	�pq�����j��=>?�a�H�+;X�Z/��j��e��q����q��	n-�l	�Uf��E��J�����{W7��ң����?S�2(k�},,2C�����/H��7C���b	HS�9a� ��2{wWg$��2�$=�i��u!���L�1$WS��R���I�ޜڍ�D�6
9է ��o�ɗ(�6Cf�C�$Ni���f��Yr��#�6���\_a�NpD���(�p�1"3�J�}�-��+_���+]�!����g�P���~&�X�z;f��&��.GQ���kat1��ކt�VAO����s��h���3�WP��n���׌?>���IH�)��5���5��J ������[�~�3IJ�G�Ŭ8D;�J�g�����7���>7���%j�Sg3�����\;�8�n�:�����9Z
atu��V]�d�5�����9D+,�5x�<2�(`��p��XLr�ne�n^�۩M��3tF#��5]4�࿷���ܑ�ˊh}0����X����o�� �ޢ#��/�V ��N0e��O+nf�Ru�K�׿oɟ31���Nt��,r竨�!��J�{n��Ir��Zx3J�|ߑ����b��@�Ilp햸�T�u���4yt}��Ӏ�^6�"��CK���P��u�?��������y���/�P��v��w���al�Ls�;�n�*�c4��FױL�W�}g�V��@�њ��W��~��ZN�R5!U�y��b��-μ��s�#8���.���R����w@�O��|����՘�pFx/T��đ]sb�L�Yb!%�f�#�T�'�nqz��Ѹ0d[�n�"��,�c�h?�U�F�� �%���a�:����R���%�aQ���ť���"x���^������F$�N�i��c��!�f*#Y�3��R�����Q ��1�-'C���_8&��Ǿ���!{Ba"F�9�e�R�Z$���Y:(�i��L=A����Όl��@U��)�]ޞ�cM�qs�)Cf�v���,�r�8�,0�G%��Aw��*NT�6�S�<D n8Af������=�B��m%��t��0��L��j������ʸ����9�#du.;N�Z ��v �0���=ǉ0����U����"�^����ӎ���|�и�Qj�ߒޤPʉ����#c�Rt��d�E��8[��ΰt,�tB��%U#.��G��F�R*�E��$�p���e'R���,@3��J�R�Ҳ3��i�;�S��x�"lƔq��I�&{c83�e˄z �\���zv��djOv��d��Tf;�� S�ۧs1�ߛ���+�a�SqB\�����";WbC�����/Ur�s-�t��Z�	�?�E��C=(�\k]4'���$���=rZ�Q�sw��:�JY�/q%�*�8#*f� ��Y�#�{3<�9����v����aE&$!.;2�'�?L�1JB���1�J�m����-ٍ�Є?q����){�g��O���gt���p��?u�TP E��&Q����D-Nr��$A;g�9˂��p�0 /��_�"��&�C� �ҍ�r"2���r��AaZ"���-cF��>˼�������d�c�x��zZ/�<��;�[n�{���:Q�:�/���Ff&w��F)3�a̳ϝ"�=��4g���Cv�R �X��#�%��@�r5��M?�o}�"	l���$�9���9��y&!۪��E/���oq1�Ѕe#>��}�k�P����h�D��x)]"���!E!�Oy�F�w��Q��Z�T<�e*J�L�ߡ����RIT�k�^	!2�oE�im��]?q\msz���DC���*2��_}��JsW��Sޢ����E�X��t�mqb�w�����MW���z�!�F�
vc���� �̕���k"&��6��[�i�u2]b�Lq�M�z�:��P9��;ɔdύJ*V?�KU�- ���&8�O�K�*V�����B/�플��סBf�N�5]g����?1e�� X��MZ��V������1��pt��j�}��x��1�!��d�'u�:�}���YZ#\Fj��9s��kz�\�*W��$6BV�x.Ƒ;%���LA&��� ��f�*�N�:�&�K�Ry���Wu�V`���l��*8V�:D[,}�1���@b؈��3�Þ�7q�#4�i���-��
,���4-˶Ex�>C2�څ�Ri��
��S�� w,w�T.]֘���+�),�ɒ+7�w�|U%��H#��B��OcD}�޹�.��q��;��@P��k�t�!P�U
j�a����_2�cj�(t���($�U�ɱ�T���
L�R�z��Y�h��\���^��	�˟�>�����3,߼Q��Tl�zF�D�� %�ʍ� ����}k+k�5��b��
�r�\E
�/�G�j��#F.�Z7k�q��7�@���.=��C�>��Fm��'��Y
}zlS4dFw����K�F��D�� �Qg�g��z�삀�cڵ�L/��5�}y��t��H�=謉���^�-�;�x9��6&|lx�b�Yk���yQd��!R��'V���_k;�_�����
W�S)�xfK���{-�q���}�̱�x�"z���A�t�j�>�5�+)I�j5M���p/lk��q�I�շ�M'ԉ'�5��;[d�FCo��iMr����$R9�	����7���I�����3!����o�pݿ�� ���S��Zv1j���u˵bԹ�b��+h�_���hr5���$]����m
��ߤ�Y��*语��»���-���=�_24r?�f�]\ݩg��x�-0���OL���pc-^��dB�zϻu��
�#B�'��N[�><��C�䟦�M��s3j���h��u�v@����|�Ɠ}�_���z���#q�o�����,x)C�S�9���`-6!=�j�&����"���E�_�������L��l�ޅ�(����n�P�m���Z�~�'��<�Rf�uEO�
ú���]	 ��C�-���~�KMQ+'��v�&ͩ(����'�rVuxQ���&�b1������r��/�� F_J2��ݲQ��o'쪇U�w�'=�5|]A`�)�S�^]��H�f�{>����a�b�`�k��
�S���]��g�9�V/�[|��e�4)3�4F-6Zh�=o�����w"'�8�U�Yo�_���IlF�p��|��"J�-�(>��+pM�;�4��*G����B?�EZ���U�|��6^��J��4���wlJ�<S������(��ZC�e�I����N��u0L�v�K��u��C�w���M���O(��?k59�sN�f�3�hOtd�t9�eܖ�����%#w̾H:���$����=c6�=�K'�ji�&$��ڜ6_R��g���'k����X�	#�?�}�q�v\���x�w(M�^�G~-f���'N��o�;��+����;�9�Xp�����QH�|g%/�}##����55O��f>���c-k׀���UG�e���*�2P�d���nA�H_�6>R�u6Q����E/;����8O��2�`�-�>��c����֤�bL܊�ٴɺ��P�B�Ta�ke�ӈk ��jSW�w~�&M�F-9�'|d��u�T���7W�~A�2P�!��w�,vaд�b��6����Pp"=���{�>�e����]a�S��X�!�Kk�����⢼�˘ũ^9'��m>���U�	�_f5��۳H��h���Q	��I��&���L)\������:�u���ï��~rF^X�Y�VdL -�^��z���N�b���XS���@_��d��0��M�q�0C�g�s�!H�OpYǐϏ�I0쮁���ȇ���E!�����n�ҎJD��G�Q=c�΅�z��n��4=k��}��E��?[�|f�ׄ���aA�Q~hz��W.e��i�Ξ� ��(�
]��"�,q��q�n�s��I&XҤ��Ȓb/$\���ጽ?�~U����nu�݀��L#$�s�Ԉ���B[�b3=�8�E�+��%Yl�tE7�/P��6�ܲ%�$��| Ed,�A�}�=sD��=9*l����J֍=��wm����"�D0�Xz^;NW�S��XX`L�v�<+B�����j�'�"��WD���>%BЦ��D&Xw8k��<���ɭ�.9&��X�=8^d�`���&I�2�M����d���1�
� ��B�߾~(^�[�zI���^
����L/Z�-bD��4c_j������13D}`G����|+Á�p���T���c�c0$W��SƑ�#Ř�3S����z.u�[��"���:Mpiyˋ�����D��(�6-}9�B�lH�x݊����c��ܥc�(�j��}�Mn�!�"�8P��^������{�_��]��Y
X6��{��{������E)�8R��<P����ȱ0��6"�d�o�Q�5���P��E$����|����F �D�>��z�x�X�,\,�Rz��E!�wB	v��*���<2huF��'���_q�}�u�,����m�4"6/ȥ!��=X���T`��LD� ���'����nӹ��VUWp6:o��Y�%���LuqP��[?4�k��r׆+���@��/O�K��?�"d�3@Q��N���r-�uz�~�%��A�ڂt�	ЅLv&�=�,��p��vä8���S��o�������
�����2�����x�_	&��Z�1rzV��t	���%�2~Z�f��������L��o�Q��y��'Z���]�W��N��	�xS�|7F]$�L�`�#��Yp1%�>l]���� #�3©L��������"eLd��V�+�MY��AP�-����[�\���l�>`�c�ɂ��[����5���T�s ���::׋�m|f^#�s�����Έ"��G����?`wY�jp��[���/��q��:��ג)E�0�����fQ�ޚzk�Jӻ�~�}7_rSA�;a`B��w?h�M8 :���a���:!��ʼ� rk�ZQ��#��!�D�;�4|��D,G��r��sCz.�P`$1�i�&�c4F�|�E%������tGܒ]�����ES�r���i��Pλ�3�/h�xJm��lԓ��r
Q����m�i����F1c{Zlҟ���W����i���b6s�0�[�/ ꇶ	��	�n�c�'Te�������Z���sZ��G q'�[k�V��aۏ���w@�XQVI~��s<�jMʩ�W}��C�����}8����d{_7&����=�VI����:K����Gmtps�1bb�ⅾWK�|�ڮ�Zk��=|5�@��[��C��t͸�Q	K7�<�iޝוgX�ocȪ�5Q���8``(2V�����}��`Z��]�Ǝ椮�s�^mhG�[��YA���#18_L]q��G�NS���:�EY�כ�Y���ۅg�}��O��'x()��}�]m�����,�%�����n�&�:�e�`3"$X����hW�̈�p��g~�Q_�ځsR��O�>Dʛr�ǳ�-�3��Ȭ�% ɮ��&�����K�Bt�e���O�w}�~^ֻ��Vͼg+�w��EW����T&ss����M%[��%�q�Ѡz��a�/q����w�ן��S�O<�X��� �����r�����A|��/Ҫ
�R�?������� 13k4��Q����,%��u����Ы&�đi�A��@3�T�>�fs�'�x~>�g�Y�:���U�\�rz4_X��ݙ�O�a`��NL�,`��d1�od�[2�r��aP)e�t�n`����!o�g���Sd�h*���:��� Ƕ+�����.�"d�R��uB��lb�#:�19\���ZnSJ?�z����G>����ŀ6U�c���=��W�Od��g�{��W��"%3�ڔ��Q���̽�_�s��Ƥz�F�\q���Q�AHI���otCɦa�"�aɿ�<�^S�0��L�jO:��}�Bx���3�V2�I����x3h�<]j�}1X���ߢ��,e�?7F�Z7���R�'����4~�i� ������A�����|U�΍�F�b�O'���4���o�N�LW���a�9��AX��É
I�s�FbY#��6��"VC�
,9���f;)�?
P)�K�$�IN}�]�8'ˎ[Wc;�� �Di_�����J*�W߇*�����͊�*�E�F]E>�̇�	��v��=̓"��W�g�ԌRh$e�,x�*U^��L_�Y%�l�������ob����� ���Vq֪���_ฐE�dԓ�� Y���H�w������b?b��iD��R�&A<�S��]3� k�����*'�m�hl1V�c��s��b����X �zĠ�YJ�}� �ñGg�Q��?�4�����O�u�U|Е�[������Jhh�4T��a!{��h=T~~�U��}�M N��������Jx����7z�����b�	A�����h��;���t4���ա]8���$F�I�:z�����{��u) �7�Fŕ���z��d�^�V
E����F'��i0]�E;b�}L�B�kzz��xtƓ� -׽���F�#��~Y���!(k(�^ޭ�� �,�WP�/����^K�ni�r�{�������=���lWc<�� \����yn�7z^� �J-��ŏ�'��,����F�z��Ƈ�Ŷu��TV�v�����.��v2&C���
Y���e��������y��2���T[�f��0�� ��(�N�<R�P`�j��蛾h��\tVlQ�����,WG��z!��*��C�ၻ�q��ϯ5�X��9]ѷ���U�fַ����I+t�|IVa|'� ����z�B?�#���ٹTz6�̾.Z+}�j��o�cS���i��x���ȋ	���������������)�^��u�.��DΠ,E�`��	IIAg�;��	8I��<�$g��x������r�i����@wIK
�"{P����������!��`[�(bбo��pkr�$��E�W���`��\m�Ԑq'���o�Ch�d�o��g��>�
[&ۜ��d�F%e�:�\�?�b�l��N:�

[��`������t������\R��^�+ue��V&��/�+��.�Q�l�	҄h��GC�E|���=�m��U9w�w>fy���<�9Hm����#$B#~7y���l� >��몋�p7e�o@�Dy>ꡆ>&�x@�em��.Nf'j9��mle�@�Dm��x�ڕPe2�qxG;5#{����%����w%�s��W�ˌ���{}Nc�qm�����b� �Z�߮��?��E�R��{�sOcZ��^��z���Q�ω�������k�R�9ٙy���/D~d����j��*T��uQ<�e���TW��io��k+2b���koQ�A;NXT��L�qډ��aܐ�F�}z��$�i�7ZZў�����iÿ~��G�}v�*�xz�� �zK�/�*��^=_��
��ڜ������o����1(��o�m���t����y>+���D��ڏ���D� 3�B���-��!��<��M	�!Ϻ��"��u��s�������a	'ޙ����u^���]�^�O��tUod�L��m/D@LBv���{�|F{�ɠ�G���3݆b�iz�BS]'�Y?�3p,7���,<�sk	�m� b~��&I0� ��S͘R��( DN5'
7"\V2ɝd}@�7&f���˄��-K�JG�ǍNk����:pJ�3N!<��/����=<�e�-�qH'_�p�"�'������5�bhe8I���n!��}[!=<��"�DC{�o�z�7�bҽA�NUp긱³����Ύː��y�0	ּ׋�'!�JG<��wP�KRB�W�͛�&[�(�I���6M%�|�Cf��߅M/��m���p/\��U���$>���k[iZ5�i�\�D>F�Ĥ����h�k~��%�v����p���ZqV�#��qL=���a,����|F�!����cwU�l�����5�I*��c���'�Q��o>dC�tP�X��)�&Ʈ� ��k� 
,7�l��6�������M9�l��o})z��lE��ѕK�]s�l��G�+�|�'��,�LJ������b�/�jQd�IVc:6�A������F����;�f�;.3q�D����eS5�.ۏ���4�G\T�&ѐ�4��e]�!�g�֩�VI���V�v�#���W~��)92/�.��a[��C��9���#����
C'���?#Mw>�M�%
R? ��%���T��B�W�ma\�ҢD�.��"Z�x��9reWCӟ"QX���:�d�P'	`��w��EBu`���F���Uk��m�]X��=b����yּ ���UC�P8q'�N��DO]k�K�f���3iN�z��C���n[NQ����8R�0a�r)t�����%q�])�v����H�16d:|�N�a��%�cR�Yi,%�O�UJ�g���h���T+���a�ɀXajM. ��nL�`x(�]`���1������(�stDe��%��sTtāz�84��h����4�ǫ�y��^���1��]vo�/�w�,8�����Ʒg)��Cu���࠲�M�^#\`nX����w�]8fXC^���e�G�5�� �񽓖�/�����`����qE�p��|Kz�~�j#�!-^�}PIm��m=�-�&�Gٗ����?A/ϼ�x�Y�����y��H[��]Pj0�V�Q�H�A9����e�1�F�����.y��J�°�Z���m�������fL��=���s��3��u�4�����Z��&��㷬\X�$��ޕ�D ]!��Eq�Nw=G6MV���jyZ����w� +���(#���&.W�S0�#T���9�V��<Nw�תD����֠-�vL��S	M�&+���7���v���h�[� a~*\���e�1������l{���9h�R�S\ZK�����Z(z��)n]�\O�'qj�����)��=4�]yu��+ܣF֘����Q��Yr��N�δ���E�N�Z���^��0��?Y����8M��A٘��.E 
�a7h�V����z��r'�w����G�/UV�,���F凅ם
bc��d�����~��e���\<!��,�����,Ҽ%���ຐ'�_3�ާ���JC����-aC�a�(c�����X=+J�AW��$R�p��+��o�H�wW#�!~xjDe�V+���E9j%f�#����Dn���U�B� 4�M�@P����f�^�RVB��{҈���(��JaS�c�Y�?��E�f)
|�~�8��2��G�.}��l�")w+b�­	�@L-&�S�3�YÝSV�E���J�F(�:�(4�,�;	��HU˂U�l��=�l�:'	�'߷^�!. �.���`o~������Q�1�6���ۅ ��-r���Y>�V���t��I#;ug#مЪ��8��z\&����n7��#��k�������L�[[9��<-O��2q�����d,�R�{����w��E6���%���[�wb���W�����P��̧hV��}�p����ɶX��:���@r��ԏ�!1/
BAG��J+�l��/����e^�\����! \�1Є���#c�g�<s����N�j'��o'�?���dk}�f�C��Ji�>4fA��"��E^��.'=Oι�F�2s�X'��Y*W)�_9Zm���\��}�%_'�L}�fǡP�1s����^��8!�+� �i���g/C�c��yP���ת1��N���C���.x�k�O��n��Π�� �u}���������W&��Tk�(��y�]ބ��
�qΖ-�n�y����c�*�AD΄������h=0����1�K���1W��
�#��"��mUV �����]\g���@:d��׍�с��΢�,��h2LH��>����l3��	� ��|H��$B�5�P[\�IKPUL�cnh�?@�������B�uH/*H8���L��B)�N�	vlm�|�������\��#BG����_N�0z6��}��؉�n��"k�$It��m���S-�4�P���WFF|Ȁ�y��z���_�b�d[�,�g� �#�g�vC�v ���=�ʎ��z��B�Zp6�ۻP�	P�c� w�݁ގ�*�AI�5��
�(��^��ycN�B,S	�<�r?"��
Q��֎���ea^�I+�(��r��g�k�p�\��ʴ:t�a������L��ݴrS�$]���!�АdT����'�����^�D^q.@�����1��{���t�ђ�$��x����f	q���{��k� Ý�>I�yc�D��:��G���|ȏ� `��혊���V����yj&e�~f���Ch�`k�7�C���Z��u�f�X��7;�z���ы"�ؓ;v�d���b�h�aV��{&�ܸS:"D�����AMf�Maʂ�Z����5#TL��X�<]�oĩ��"Qh�xsc���+���'K�q�id&��d��Tn�j�uW�\"��죝��0�C1<cC0sd�'7r�h0�-K�DxBiZ}|Gk�ڊ�5*埍~�b���XeάP���sk�ʼ�B������rgT�<�1���q�U��!VvQF}���CBc���L!����,uD*|鎖1\3=�VkD�2'��AQ���.�}}{�,��/x&jid�n�.�Y�☹�rȿ(�ã��	��
���8����n�&׮z�Nۀ���C<�r�J$�5�6
La}
��t~��#G9J<B��O�:�)����  � ����գ��̞/��(רq4~��)WD���ێ�6���F:A��\��$fwCz�cB�"��5)g:3�Z~��({b��Ϸ}�1����} ec�����zD�A~��U.p��X<Tnɲj��9�/ZfN5>ZPw�`�[�Ӹ�B�a���"��1i���>J�ir'Ԁљ�g�Oty��*�3�0�i�M�Z=r��?�� �{�,�����8��~Iݗ��\�3)V�v4���K���!uʅv�>�i�Ԙ�ٶ%�8�X���8����9;ɝd����	�lA�ښ��1dq��ᑾ1F�0�����"�������l�q/��:���M�!a�3bI�b�9��R�?��8ĉ�13�:�ـ��s�b��r��j��cV��覢x)�jb�d�6��j�r�_u"��[_-bS�C���7ψ׆����7�0c���,�u)�o�⨢�����`QZ���+7���t
��7*�U�	��'t��%%^U������v\�6+m��pk��O��<$�mMl�����ўd�z�����q�c����Ӝߞ#��%��[�r���x���j\dD㔄M�t�	��D���Z��Fû�1�S��D�t�5I�dq�0`��p�M�a}ȃz+I��xX�+q�pG�[�_��Z�i_Ӻo��H<��������"��L
3�H��)�(�3��-�.~�E�fT�/��+ɫ��ӗ��������������I_`����@x0%t8�ȣ�OO�^#�ᨣ�D�k��u�Ʌ�hM��'Q�E��K3�$B�H`T�䊹0� {iGF �G|��?Y�5i�MDc�[�F�	��~��� *�:g H�d��j[�ˢ,���~� P�;���@�;�ҁ�(><[z7qV0����j|�c8۬S�A�,��(f���6�4��{��M���j ����@n%�k"hװYn:d�� �X���la�Rs7
��0,�(^�F�����'�h�э~w�� 9�K���i)(�c��"@��ԯd�3^"}����R��V�+6B����']���FL$���·��7%�B�8J@��{f��1NG��D��%J�	����Fz�����*�M➑a�������r��j)�/��^zO&���&�Y`�|χ��6����!�Z�x�bo��4���yj�
<ZA]IO��=[���u�52g�@ ������틍���N�K�����rD7�����+{�Ñܤ3���L��l(���I6#����#=�U��V��"�e��`�i���т1�K�E�z�J'�P2���i~�P�(��)'Z�{Q�,;D��|5)*9����Q����3���-t��̇���ٗ������e�M��wd.&�,zw�Fr�K�ߍ$I���@0�؏���%(
���:�J�\SHC�	���_Y��J0aXi �ϰ\���]0u><�n�GO6�r�t;����B����G�q~���`�a��i�'�nJ�k������AH���Q�`��t,���M6%��8d���f�,{+ͻN���u!{=~�<��e/=�5"�:a�FV�Y�ҟK\�& ��f��]����;�����ρ�5�}�x͙"#�b�#�jB�9��W�-��Nj_}v�����#OY�&p\R�G�bL��[��i�yLۗ'�53lܘ޸-�e<�uB����MG�j��d5�n��׷�	5[k�Y씼�zN\H%�D���{��5�b~��$�{�4�` �b2r�s�� #�Ik�/���q"��}�(�m����f9��Y��s
;��~����:��@���4ܖi;I��f2c T>K�6��+�ab����s
��1�X ��'N"z��~�ȁA�h~��X�g�w� ����^Z���E(�D��ʊ�i����Li�U�k5P���ߤe��Fu��W�>o�;3R��f
i�Ofə��P����2Y�FB���C��C�S�
h��L�]�B�E�7�;5��5��
���ۊ5	R�R���aP��+M��%���#�x� ���¢6�|4I��ױ.�.v��D'�bܓ�� v�f����g'�I�0� |�L3�D�fvGN�#�s*nBS��p�xP:���Mp~#+���.�π���/��w犳�2����G��6��RxE<�6H���D`:��Ѻ�V&��t�����AM�9�0���]�Ι��~�R�S�G��6�	�#�0/!�4�n{θ�1��_��E�(���j[#�P!^i���3�T��J `����ڎ�g���(w�#�fzcọőɼ�|��ʔ��X�;�9�դ��)H�;�y��{9�Q�_m����zI�P�|��׼R�E��Q�0jW����*���*ǁ�5�F��C&I��h!��:D:���`s걆P�������.���f7=�M�?we�:U
������%��[���7o)��7Y�#9<@3�Ç�#���� �!8��֨oms���K��WV4����9��_��X�E�u2����6/ً���p�=i,�q�]X)Ę.�i��d��陧�{�����.^���5#��U���6s1�������d�N��i�|İضɼ���n2?��i�H�t�~��,�8����hwTE���b�������L�c߀*k�./�RH�!��}��a+�spL@J?۽�����{T���=�̺&�a�	�����9곤8�V�~޾�����:����\���N��f�n��Vw�,(���S7v�,\��-*O�r`yU�A	�+����W𿄌n����f�%f��D�8��rG�5�f.S��S��W-u�W�P$L}�/�wTqk]c�Q�,����K�\���g`S�gve��/d�T)Sx��?���V����mT��k���қ 6�kO��i��.B��Y��C&NK&tu��dM��I3�D��I�OF��`B`rp�������\�$J��_Ȣ�������C4O��ٿK���%/K- �)� ��^%�-�k�6���XF�+�ul��e��'�Q/�A_F��ܹ��|B%���$�/�<�Pf���Y4n���x	��ϳ�Q_��ufUr���W��ٴ�X����Du�2w1Pi��P�D����/aUc�E3g����wg� `	��$�a�j��m�\�%�|���:h�Ǯ�|q(X2m�Jd5�� (�f������=v��Ҽ��؋��׷]�{W7Y�$�����1t��Ie&&p_��)���O.@;�7��E��)g��^=Z��^¨٢G��<$�_��a'%�fLne=!�m���w��}�K1��tKK�v��3B[ض��u�8��wen@X�ka;�F��2cE��Q���ix�ߒNf��D���dA1U��OKp�\��<��4+a���mʭ%]z�
���+���P�:t�T$B1���]43�-��&�NmZ���#��H'*&���;ht/S����]�c~N�pAp��5)��� �A�A����yO����
b���K�
�r���c�:v��=�@6�9)�^Z���6��Aܙ�ut�(�kp�����ki�� τ�fh?>�����'i���|��Y��4�6f��⎠���k!d���Ko(��?��c`dY�q2�'*��6��cE�@$N�{X7����&�{�T��w��;���r%'��O<O�X'}����o��uB���(rB�ei��"��2� s﷪��jC5�^i#�r�f�a����*}ܣw�{��������86��93�,����2���|�b���ʒ�`�u�",;7w)|,v�zF�;�/�����:��}�������z�N�!�T�9�5���e[��7Ɓ�L�~{�}1�D��+���tBr�J� H����ȉ�`�M��K�p���~�p�t�p�L����"���v���#E�������X��@:�U`�o��g}%XcSӧ��)_a����d[�9�dȷ
_��&���Σv�Vqf;Q��1\����6?NW���J���i��:M��g>a@�-�4���Tx��#%)]���#�o��ö
KC��b���݉_P���u�uT���F
+��ʑD���<r*�E8��5oHg�S3��OO�f+[c��,V��OٱD1�L[�m{^m��{5Z&�;��$�96�N����H���hAB�v���ʅ��ِ�����,g���B�������x���P��e��W<�V��IN<O*�-�iu8$*O/�����ڤ�' �D
����&��n��`�j��^5c�nZ� ����D��e���h=��г�?��F�021T��"�G�'��:�6���nq�v�uIB���m oD��@���9e*�Q�'�f���v_Ո�`W�f�mI����ڹ�1�ʥW��UW0�)4R�d,�uOT�����8���� U'�.<��Ϭ�qY��m��3,-o}�i_4�?`���ِ�I��^[��g¹���z^q$=KɝŦ��/�C[�$r6�3�9h��Y��h����T-��-�躪�nh�Жi3A�+Q�ʘ�3^Q`|�mcF�qXF���,�9(s{�j!}�n��Vh%Z�y�A��n�1�ףIIY�DK@��z"�����]i<e=(�[����H�1�P�-��`ͅ��!"����mϞJ������+7~8c:Ms�	=r�.�������da���^�	e�Noc�"	���-ɫ.�CF���,��̺K%F�&�7ĵ��:-iW��Qp�0���=?x�g	 ����AT�a�\��� �ъ��q�z-��*Ĩ�k� ����G��/y������@d�f@��%��p���{�����R���g����Fз�^��mf^ۇ��ʆ7B�Qx_����#����	�'�I?-�l��VI����AS���@�x	tFo��Jhk�q�5�엉@�<�9��뷳����ⅦNj��C՝�/�5��g���;����H��x���R퍧�h���92Z���R@3p�m��ۦy۴�]�*r���ͳ�F֟k�M*�$��׉c�qA�(��|!,�ad0�Ѱ?0+8�)��	���,k��������B�U���=~�s��Md��k9w�$��b�̪@p��>�<�q�����pπ�rSg$�uuA���a�6L.�iM�� y8�X�ba����6+E�z����m��7 ��}��.�H|�������n���Xa)7���P3>oζ��ou����I��q^^z���|=:�Ŝ�ƄF�e<�{E�d�2d,�T- ����=�4�"גۜ��YrWB߀]}'n;�	�G�B�p��+,��������� >��ȍ�f�������h�S���!L��&(-G�<x)9_o�K�b�@��5�~9+�0s|[�����*��M�̴�4��������Z�ys;�($E'mf1�6��]-�Ƶ8ގ���Y渞�OHx���=�-�E��wD�<���9�?N�Ym�},u\I�e���9�s�]���[�;iM��@���~Z&����E�	�j�[<��nb�ͭ�R�����"]��L����Ã�#Vlr���l7i����R^��x\积a����*�e��d�Y1r�O������'$G|-����w�zU!��~�{�p�.+P6�y
'����D�|�"h�-���ȝ/�[K)@��;�i��w�V�~ߦ�~�#{�W�ӓ�h��vb�M&���{�h�|�����~�zJ�Zh��\�W'�q��t-\ �9�>��F�	��ƟN��;<3j�@�Q~�S�$k]��\��y2��Y�8��R�n��;�S��O++�C��!{�~��A��w>��ej1[��w[IӗRb�h�<|�������Vţp�m�h�u�:|/�x ٵtw'�.Z�����u� )1Ot���ٺ30腼�j��{����藩Z0�/N���^�F��ܤ�r?&Xm�E(:���X��,z�2o�כ?����O���V�R�h�Dj�a���^Z�:][�
՜|�Fr��~u�9RI��R��]��Q��������Ezļ{��p��g�\a:�.꘹K�|�l�|�p��P.�K�R����G�X�x���dZ\�y* �B�#{]����!n_����=��1bu\HZ��T[s�lv.�8hyA�=�����N�= �Z�>�M��a�F#�A�ϲ��s�������7��IqǋRHn����c\D�N�K� g�1f?bX�Ȗ��!]u��r���;�"�-cOS~|��<*����X#���b������o]&��n� |a�6�lǧ������ދ���4ۙĉ0�	��q��W�Vp�"C�j�x7�cl�G�Q�3��9��0y��bPǅ��#T)��#�:������Qs�]A[n�|��qx�C3��#��2>��DI�V��-܂�(nYt�uT���_���1���үb�ܙ��'�H����#g��yů׾tՋh,�S�����Ũ�һ�\X�s��c���ֈ�<��zd.Z��1�Y��y��� ���v��z�n�,������,��W�@�,�>�����е��/+a*�R@��r��
I��*�󞁟{Vۚ2	�Q�ü�� �������9���ؔ8�=�Ց�cug�6�:O��K��*b`  0��X3���x�	}�q�c,?$
z��ā�a�	A	n����Z͏N� \A�@� �)ţ��fƕ5�����W�"r�uݲ���er*d�<�!�����|Be
B�ޟ>�ByPUiK$��MԦ�,�%B:_��"_��
:��D	��qg����9��/M�N�8�@���/�8q܉߭B�&p�l#��7�5O�4R8�[+�5_�Ed�@x������.��d��R`��j���b�p���`Io�	%�*����)%�nP�a����ntxK��E%�:�����wM	_�����x����'HȖ��ۈ����!
U��E%+\S�#2[Io^n�_��]��Y5:��f�v�h��V~��۔FΊow�=�8$�����@-]��`���e�E�Q�a9yg<(�͚��v�Y��k5�qb�K���G0��Ln'EH��B�?����)�Fw���"$)�_Ճ�����1������4Գg4��eS�_�qa��KU�e{�HQ��vz�xڏ���Z0-�w��� �w�}���7�bЊ+0rX�F
:�Y��0�+�Eu�K��E̒�>��0�`?E�_���ީD��.T��i#)G���V�s���׊⽴�}�)��%F�l��w?�Xn~P�pêG�z�^-�N
�\��(żݓȑoѓ_�wq,`���x���/�Ng��E �:$Pd�U]��T���JYo�zS,Pz��;:����-�0��4�M:����2w���S���/)��^���:,�C��8�(>
屢Cm�g����Zk3F�jQAv�K~��PWa$�Ͽ 5�G�̹�p֗�}apH�Y�)�?m�%-r-���%��4�_�b^t����N��_���M%�ژf�}�u/�n[BJpâ�k��j�Gȡ�^o�K�{�Z4��F*�EH��$�����j�Wp��=��D�v�@u��UX�v�Gzv9X߀0R	_���H�p�����ʅr^�� Ǖ��s��QI����/8��"X�1Е�r�w<���B�;M�b�U/*�A'/�'Ĺ*6X~wֿ*�iV�hwQ��&�Wޡ�|ݿ��2D�E
kj�P��4`��\pb�5�qIi�Z����L.�
e��6!���A���5��-��^�s�~U�޸��[r|�+w
 V�H�N& ����*)@�{3P�����1�F�۴}a�dqK}
����l
>�=֦\�AN_�O��3=���^b��w�,dY2E� cO�U�����I�W$:�n�օUw��8 Q�}#�Y��rх(�Ȳ��m�2 ���V���L���-��)���5B���sʡ뜴�����oW�i�˭�V$Ȕv�t���ICp_��yb���_�jY��M���//ﶤ���������p�1��`}�������`)a�׀��К�=���\Ϳ�w��l���vq܋A���k?���"b��@	f�r-���#�A��#W���i����2�`s���W/
�|�a�!���~"����@�C�M��<��`��Đs�5�����i�AMY�ⵉ�v�l���9g�l�i��~y���F�5󠦿^ϴ`�L�L+� WnB�߇�ͭ8ٱ/�o����>,/�
dG���b�i\[�%q;�}���Xh���ݘ��T����d�6]c�FH�1I�Ԙ"y9�t-��dx�.цr�*^��<�p�ɩ��M�؃�6;%G	t�ِ||�gc1e�u5�8`��;�P���'-���K�_�)��iFV_&���@o=��C� y�7;Z
��L����4C��$g��<�}6T�EwX:��qv�X
:"^�s=v��W��mG�zԊ���U�"u�7�5���w��0�?�ugX�5�G������]��G�Rx//�k�z��A��w[}��|��-��*�p�����=�Ab�^H1� ?�)�
8!V6���οTʭC��|j�.�zC7�$���I����0Ҁ&�2��]��6%5�`BY8[;ʡqݐ����@w!�w��/�!�^u�$���5�1����usʄ1	�P�ʬ�\�&�N�ى��)����#�A;���6�R~O0�ioF6���d�phI"���z�2E�x����D��c�Ӟ �x���I.Y�L��v ����wNH������K�w ��c�L�Y�f��*����2���t�-I��� U���e~���d� �����i����� ���R*}@�Y�����DA��X4��Jb�[���	ЂM~u�~�H/.�c�r1C�ׯ}��q��E�=
r�X���������U�>�8��8���X�y�K���s������������!�;U#~�άl㐰�N�*��Ia+1�#��p|γ�������lLO���P.�&�@l�&_���Z�������U�Hi�d�q�~>NYξ4�Tߣ��^�,�6�pԿtw������˚[I��y����՚���@����ݭ'����}�F�oE�䤚F#N���"�JG�l ���6���|�:�5�%h��(Ԛ3���=�:��v��{[��/O�-wb��1��j��e�ͺ
)�A�(}��>���	�7&A�bx[�Uڗ7JV�KƉ�_^C��s����<x�ɋ,Q[q�X2�5'�y�V��X��)�s>u9'G�S{���!�]"�R�z���Ds��zr��:�圻��4���n�]��ʑ�מ;�r��4 �`A�J�tU?h��={rxe�� .?1��P ���`U�����Z��.|�\��r�鏈^���Q�Ȣ_���q�Ҍ�$ּ���O0v�)��.^#šI$�:�P����9�B�ہ�h�Pe�A�9�+L��(�@�k�6����EO�]ۏ�f	>g
\��}�o����PZ����S���$۽rC��n�+�b|�;�2n=F)�&zb{�v$�h��`{N��	��0�ɟ�&D�D,DLs}�a���l*Rڔ�pyO��|L�ߞi%l�N����O`lV�8k
/v;��{�r�����_���.�JgV$�^��r��|�SX,���o�A*`�ɡT�g��/ci���m�8�s>"|��;r�~wIzi�����Jż��S"�MP �th��J�̲<P2��4L,U]�;\�k1�4컧���ݵev����8��8�Q=�����o��ݞHUM��O���+ߜ-�ιBC�䝽��T�9�*�5�����z�C|Qd9Ȇ��E�D}Jx��ܞ0NYo^1����ӕ��ZF����j��W���MD)�?v���;u.k)�v�$���4N�b�u���Ic�(��z��}����s3?pٮ.w��`m�x>��iyT4MˏyOW��k��s���1g�a��kNVls,	�UC�F��5����U�fbtjA!P��-h~OSv�68�.�Z�t�
�B2+%�`�.d�A�\�4}eX���ួ>t1�R�#mqls-6��n���Oк�\�{l㒮S%�F��Į,Gq�PÝ�B i��2�֮�Γ��^ؿ�0Jj1��U�~�7ew�y�������`�b���QY�p*�I����`0���f�T~q�U�Nq��n��Zŭ�,NY�@�=}�RHÚX���'�����.�A�0n�Bzld)lh��G!4֜9G`��x&+y��9Om�z�<������K,��:V����p�͢
����@}����ٓ0j3�# �픂��%�gb�u��ο�ܽ��]��>�Nz��k�\(t��}�N�'H%��z�~�F���j����_����~�a��$�JL�k¥K*��Z��I��Lݴ�bP�P�:����lD��"Fٺj�u�Q|x���j<.=W�a��(L+3].!���\��"�J���+ϑ)8L�y�(ي+�a<$T����6!��f=����v��JuS��:��!i��Bv�ᨖ`�����X���?1Pw�J�z�|۳��+��\�C�-�!��º?c�q��p#U/>��7,��!��k-���p[�ꓟ�`�'�<w�H|�n�1
��pWL��}��)4m��9��c�xr̅b=��`�&P��y���f�.M�7O��K��]b~c3�8��Z�I\<0�,�����^�Z*�u��.$n�D���0NB���![S93�&�,�
��kլ�b8�Xc��Mq���ʓ�F�� �ae�G��C���z��n�<��b	PmNKX�o�E��tл0�����j��L��Jo�d�k�F����8����%�Ps�B%(u�tG�ȸ��~Y�T^Cm�ANV�����V�����k,;!j!(E=��0�5%�V,dؐl���5�o��mo��u�I����6����3Y\D�F�2�a����$�����v \����bKz�K�j�w���L@U2�e;aȵ�L�S�m���
brY[�_�?�P�?Кᜒp/�'����[����O.%%ғ��l-�	VN������ts�Y�+�$�;�M��uO�	��%����������������9�
S<���N�N��VIh���h���7<	@Tܦ��O�����2ʘ���ݵ۫����?�"�(P��$����؈�k?J3��V��N� ��E�['G����3�oc��ƽ����k��#T�Wdۛ��/ELiˇ��R��h�0�{>����0M��)W�&����D���*\-���w���/e�&�<��:׬�?j��XL�$)���%r�Y�a8���J�!��Q*�?��֤0��$e����c��h�������;�Q��;Y	b]����8�c�h���� ֞=Sl5�$>��g�Ż�m4��/�l�S
��%qW��纊q�=�򺊛:���i�mc�w��u!2��6,�[ײ�{&��h�/Q�D�b_��M����
�=_�o��mP��R��w\�-1�I35�(���2o���GvӍч�-uco���ͳ���I'��Y��M�@d2:a�ǉ~�nnX�5�@-8�*��\�0;�5����-�/�����<n�]��<���/��P�o&����+�ń�g�·��Բ�� z��U�Fvyop��or���X�I��fӑjo�'7��O�&����C��*��朗�^SrD:ټ���^�6�4&��ɁoSڙX]ɰŠ��2�5k�Ŧ�����@���@bc1@��@@��M�05������:��?�^����[�����x] �"ߞ�t{�.ь�y�mB�DpJ^_R���z+�l��:9Dk��Pl�D%��1�n]�l��AIJJ��춞� ���S�������ЈB��q���>�LK:�d�	 �*��ۀ1��o���'�J
�����ʻ�V��k�Cj�A�7_��di�4���U1n�����j���.�js��X��c�'�v5c�� %l/�?՘Pb�s;m�C��{Cp��JP���L�N��ǔqF�G���a8��BB�Uim�|��&:�9�}�v����Cf1�������B����Ȉ���M�g�� C���Oi	���ԋ���L�£F�?��Y��Q&t<LԱ�il�����!��nK��T�&ԔU��	E�`��o�T�x�
l�e�ICy�#O�-M�$6�ì����^�� ��i�ַ�<��P���>�>��i^��~6J�G,�
HL��kP��w���̾��ojn����p�Qz!�=L�q�B�/�mC·�j�����)�.)9�xD�a��"S�E�?�tG;ћ=�ޟZ�V�ɡ�ܮ){��x9w����#v2�mz&�a5Fs��=�5W�[�_��S>$�	�/�R�T6���<ڧzj�����)�2�[�0��gA��A�<�V�����Շ=������I�ͣ%��-��/�$Y؀�e@ۣ��O�����30˝�q\v++���R���L����(�ka����"��_$'=��QЕ�Q����3�mI�y��ty���hq��[�:��@�n)���c�KL�j��Ա�xl;��@B ���FN'���kqJ^d�S'^W8(7�i9�`�b0|���'cƇ�E��r YfN���+�d'7;��%ip�d2w����.mR�^�F��jz�'��!�����t~֔�J�B�k��^8����<_M"���F����֓j����)��p���U@t�]B�n(`�_�*9�W��G��,@P]�(m��y�)V�y_Jȵ�j��5+м ���O� ��v���Y6�ߠ�=�p��V)D�^*k��������1�gR�.6�1�Y�V�j���숪jI��B@K�)���ΜWI�-|�4%. ���(8�	f���b��F��_�(����pC!��`���$	W���I�$�js&��"��ȇ��\��99��X�U�,܄Xaء9|W�ox�m!wd��)h�0ء�YΧFi/�ȷW��ݣfW�`�P2�6� ���<��B�b�oM��b�+g�t��lI�W�8�O�뻐d��H�f$�0�^���y	9�''�\�t��$m2�������"vE������	茋d�ʆy�y��˸��őJ�$B��&��Ά�& 0V������|�Ws��R7�̂��@�dѩ��Ռn_X�Ӝx��TS'��yu@e���$L	ZW�]���F�|5�J~�G�vh|���F�5�*䔙EHsB}��W�jZ�4:�Q5
Ͼ�ů0���p�.ZY�$��$y5އ{d�em��U��iS��*G��M�z�D��G*է��VQS9�>f�R����qҌ},�7YL��p���|��c�gMm;e�9��̾"����x�E'%�p  R�|��{��Z"�Ym�����IW���. � @�6�"�������C�Tͥ�J�I{5�����B�����mf7�5`��z6k땞/ǡ�Ք��F���5���;��/9A �"�^2Ӈ7�(T���1H�J�����t��˺�m°/X<T�K��i-ϸ7�{�i
|t���6X&��-ϵ��{��l̛�t�y��(��ѵ-���갂*|��H��y �f8��霑�l����� ����F����U��д.���ON����z%V,�%�WB<RU�~�/9{�~E"�H�b#`1MY�m��=�>��r|nf�C��y ��ɀ���N���2��#����m���j<�ǿ4����b��"U9dF��\m���{�)6�2=z|��:�
O�1���\7ir���C0ݯ�g{���h��LB���H_��Qz݆9y���[�ȥH7���tWǍ��a�۵ʨM�$\�J���gx����E)q��m�T��W�9�����
�W���w��ĕv��V�'��i���F�=f�R<<���9}�r�% ����o¯F���#�#�n��䶂���}��F�n#[� ?���2��-�>L��򃸜_�GR�Ff�������u~����Q@5�%|�P���	�joct$�7�$\�Zo�7�L-Z�!�qz��CB��n� 	4[��lJ{��U��D(C��b�m��b��_�8�!E�����͋�����b��m@�h�Ħ�B|�wr��'�"�����O�S��U��pGkz��	t�GM��tREF�䇝*�'�����)D���t�R��f�67�j^�h-��^�>5��:��ξ�K"��+m�Lr�-\l�����zM��(�c��$L�_	�K�0��m�E=�G���*HĒ��&��Ĵ�[If�/*ښ� ��q��k#0ʰkG��0}���k�	��1ƃ��6h	�!�)o�����(� g��h����d�;RG�7 #�C�!y?v��@z:Kj��)F.��$��9*��Qe�`O�SO~Xz(K�����ɕ/���L>����=,�u���+����T3�?��S֕�?ůLLֲ��4��H<�ޜY>�hze��l�h�)��Y�� ,����1���o�X��:�W􁇢N��#���c+��*�H��,ʁo���`f�d�V9��R�����
D�ݬiAk�z��z�c���!���KH�� r���r�^��6!%D������4aoq��r�|�n�+n�kVYѷzm�T�N~�C�*Z�>ׂk��S�зǡ:L�K'��z�\��sתWrvi2c!��@2/Ɇ0���	�l�����Ը��N�qݳ:�#dc�BeNG�H,B�oȁ����N����p?k�B��e�D�j��ao�h��|�v˓?�o"�N٥d��;�"�*Hg�9�{g�U��,D&ͯ\����G&*��XkdD�m�nEK���8@�Mo��D��$Gc�7Q�8�v�ވ��i���^����Q]���%P���:����m��K���)0r�;ڎ6�XA����İ���n��_��Q
�������?x��vLe�G%�r�t:B��"�H+SM�Z�e�gp�گ{�9�Q9��+�
"��^�n}�Z1�,j
�߶3�V�#{G5K�S����aQ������5���u��d����T[�B�5�ų�ܶvE�Iw q~Y�n���}ƇV37��E=�ݴ^��Hoe�3X��xq�N��^C����,�1�aK��[F��t�0��tz�ؒ.��>4�K��d��Y��z���#} @�'��O�э���EKdgt؋(�0����Ɗl�+�~��2�?��T�N�Ր�v9F�bm�#���_��yK��P?*
u�_qv���X:�/*XdmR����GcL1Q��􊾋�ݘ���e"9��H$�xI��jq)��r���x�t:`��s��E\���:��y��oę�ᡲ	Du������̫c�?�jŋ��ksr��==�r¤���L��QSy�%�ǧ�2�-��j�6�ֹ��u�����V�O[��-\�ϑ���K��B,'�\�;ڜ�``�W6��ct�$Uk�"s-���+����no2�����!����?��|�9H�e���q�Jv����S-�)�����X���������2�����kË����v�]{ɓ�<n�1�2��Гr�y������VY����4E�Rm��5�ɾ�Ҡ�)�����\�݁��5�B�WŌ$�hxB��ؑx�S�G�J>���U;JQ	]=+ul���J�|Y��+x�״ؑ��"��
9s�y�~� �����ŏ�ꑀ�'I.YW�y�}��f�W��!ζNR�S�D�#oLV��I��B�jX/�(*|%�����巀)3!L�P[��O��ln�����6���YѡT�a]�AS��:u�:�����=�Y���.A�m�9vA��S�N�Ӄ�豤.�Ӊj�4�2��^�|U����oe+���};��+I�?���8�h�-ӧ��U"���`�밂����`��5�L%�D�
�q��q�n"q�3}c*�G+%��p��~N����D��e8)�e�A�� ��Is����t�zߍ����_�y�������H;L�cQA�6�s���|�p���@j���BG�RB��.��81#����!E�,l�&N��Q��$I���' ���[g�:��MNmVTWi�q�o���>@�b��&����7��E|�<F�۹����$�#�#��c�f�W �1�"a��	��dK��c344�/�g1�)���Ȍ�	&�J�G��Gbd[2@�'K����:H�Pr��ICr��ǉͧ�B��0�.�|s
_`&�Zn�.KqH�,�A���kr�����S��@��k��^F�i�458�P]'����.���,���g)K�m��ՊI�ҟ�0� ���p5x��Z>'>�� �(<���.��h�4�-�0Y�(�<��k1�:�2� ��n*9���<D0���,�H+�*y�<EMƢ�%L,���-}��C��!�l�6Y��x�=��%[���H45`ZՉ
�����҅z���B�sL�e��}a��Ko@�2\�*��5H�v:�D���1s﷥�h���7�Ȯ���׼f�KAF;�-~��l��S� ��Q��V%��%N��i,��F9c��C�({E7��:�U3��.�B/���}�I��Ylz��� 9�Fa-d�������w��:� �q$�ϊ�%$܄�Wh�[���+`D�tH�*=X��%ء��;��	�L��<���W�Ei��'h���>����Y�7rvk&�a�;;�����qx$�X�:q��6;9L�^�_�P�
ي���i�A�!AJ�@�e�Q.`�s���6���z^��>���/C�ˍ�Xs�9��쏇<A/�����(o��N��5F0���E���v|jW� S�oM�d\�+���h������(�b��F�-�����e/N�a	5s9�-�5
_������,�԰����$o�p�o�����Y�g�G���Y��-;���#P� JZ���c<p���rM�T�]`� .7���{]4���i�wS@ �ڄ�^�ds��3?z�o}#��8�i�����+07'M�j�?{�
zٛu4��(�7�Oa��}�*���+4*)��i�*j5�Ꭹ�f�É��l�g�a�8�H������{��高�b�5���\��4��):d<�u�5��v,��nL���;�*�+��(�?]�tLƈ�Q0���O�i~��F�,^�ۚ�>��_--�t�����E�^
c��fV"���נ��_���?�lqvK�;��Da��(aL�Z��fy�P��{��s`ڲd��k���v�n#ו<�`3W��3��5�Z��U�<��Ӧ�B2������E��Z�zP��֛�����0
�+���<3�T�π�����4�f���Owl�!t���s0�����P4��/�D��g����g�\VT����~���5�,�jg�Me>L����Za�2luB�~��
c`]1�Ӽ��㣶Y��.#~��ֲ�')��v�����۩��VH�G�2G`̻{���䢵��l��+u箐���Јg����SFb�������8
0�Dd�t��T�����*�@$Z�����/��w��&CH�� � �J*�Ãў�MU�E�y���$��ÒR��r�#8���b�܏R	��BՕ��LN�[IFv�p���E��/r��`$B���~Ѕ{�^���s��?W1b�ӣ��R@9Fܥ{�t�~fNz��owX����"�~���p��[<Wh��%��u���q�*���`5��A����n���$����`�\9)HUדk�s�-�N�x�4}�$��.���u�+����k���wT�'c��#
ƾ�a`]�T
)�s24t���01���{���6+�O��S���T�Z���y�Y򖠘Y'f@�Z^���}��O��{�S@���l$`�&����o���C'&�:�Ȓ�C�S���D�����T-dWH_�IN�+��o�G(0��Ġwf�Q��f�� �#(����c�ڼh����Z�-O_������TQ�-耴kC��8�>~�YP>g�)à`0tg�u_� J��s�?����o5ID^��ҫz��[�����Nv�����5��\,���?����!Yܧ)R���ΏEJ�����E�_���\٢J�>����/�)80]�[ן��o`�E�U<dABW��P�H~����J�����u����hH{��@�3ֈ��k�c^8��m��k��sr���+~����=���ݗflk�pZ�������Jf?~h^��H'�쁩z��8�"��#��ޑ�5[��}��w�G�_bC˽�-��`���D#P���3T����]�K��o�#�Ne���/y��`���q��-˰����B<;�K������v:����3w9$��?�y5�`X�կ��T�}NJՁ�b.�`(�mJe����	� ��D��:B/����X� ��m(�����t�^[��s=����gp1��̹/�P��L�o�6v�����I�.v��4$�>@^C�L����6���)+9��Qh k8��d`Z!�boɸP�<�46�9q5`�"*X������"��QT-�V��%���%�U�7���Dq&��	��/��k��d���
C�% �l��"�Z0��h��d�w��u<s�h�	�Tp��&��o���@=A"�����S�Ģ�ݐ��#.�G�+x��(�Q����#k�+�^��툦$f
.��Yε���1�bU��2��1�Rr�/|p�t^���!aBkS&� ��U �:��B��X��x�}*ۥ�,1���A�4�Z��vE!��|��Oê���]�\����4M��Ws���$��r���$�j߰���mhU�2�<��������Yi�"�����Z_��~.����[��4F�WɆ0y� ]u�6{Rz	A���� ��6��vo�6�����c�����8%����J锑A��`�;}g᠁���9����W��׫3��h`�q)ys�I窉�;FɆv�l�`�-Xe�Y"2a�O)����ؾ�ޑ��y���7��ɓk8��9�O�v�|5Ot��ݛ�"P��⦊V�b� ���~܀׋b��#>K��.#ҴL�`b�@ {Qs�z�)�olx`
������3�x��.�@ <�Յ��$˱g<e�"E����m�X���:/mo&���U-m��\6�F���C�Rr�����WЂ���b�4OkŰ��ݔj�l���L�q?�;v�����n�~�˜�K���j���b�F�U�(�d*C�
Q�c�#���9�9�yV���_�vLp ���Z����p����zO����`:g�6��)Lhrd�GmE�C%�ܲ3J+��8z�~'_|SڗMQ����| �9���ζ3L![��3sT�@T���Xg�Q?��d���Y�!��\���M$���%�>�a[
�8y����U�B��`_��KLU5���Ģ1�	��R��qR�����0�%�L#᷏����n?Bg@{�>>�m�ጜ�҉�7�;�ζ� �C�{�)���ol����6����V�w��M�� U�8�.B@���;N5eHB�wv����I�쮵�Й��\������_}lZ���-+�+��K������.f�RINo��nr��g�)sE�ht\P޾b�}[cuc�RG�J	Px(ǒ~F�7�H�z5��"��MWC>�[���U5A�[�W��t������w@��Pϡ�%B�)��/� ˸E[�huƑ��>�?/��5���1KXO�R�'�e����ҭ��V|P?���M��}�ހQw������;E� �}�o��ۇ��O1�zSa�sKx�7����2����uyް�O0�‱��������zx��{Gz�z;��8a�&}��x������d.I�>�@(�~-�	J��������v�HƬC�!];�3Q��a@?r2#��!R�6������k5�o���A�āجNn~'���Z�#d���*�݃���.gч��[�JtB�B5��s-x{7�2��	1z��є��~��k��g�%]��C��`շ�U�OV�gT9N�U1x�5��7㣸#�䒷�c���knΖ����Q$l�ď)c��)'֋d�|rGu��8n��J���O�ќJ�[}=���3�7��-a�?��d�hvk�5ś��������c�F>��!dz�aW?co�<����BNb�@VK�����q7#J�bXn)Fp@�!�I1mT5����|@�؂R/�����HX:�O�)Q���><8F���M�y�H�Z��Gߜߵ�@��?�x���\GDa,z\ؐ赘�� ]0�v8��ҍ,���f�8ѯ�������a��EJ
K����W��*���=x�+�Fɣ���S�:��'=4�o6'm׊q�F9(�J�e�7����v�T0�Q��t�?D�5|��c=��fp���Q�����{��>�`D)?�T}�f?8��.�/s���V���kr��@�,�?��](���D�ӣwt� � �<5b���ӫ��Ƨ�Q�R4��a@i�B�����AT���1'�!�=+�%�9=�v��@����F�]�NZ?$k�%�zhE/�~�j��M�±��Г�sa<��U���H�R2�ȫ~!"6�����$E����B�5�ڲ{�u�ry�( P�y��6"#
�Y��_NdsFZ؎pj�eG��|3U�O��\��������:��*�與��i�K���0{�@|�Г	�o�e���߬ȋ{E�xׄ�J�y���ڰꞔ.��m�ڟ���E��O�J9�n:�� 9�=b��H�h�۫�d��99�1�A?0����� ��+� �R�T���)IZUF��WT�n��?S��U�'���q�!� 3amv��@��OeA��~�DCE{o�)��e�y𻧩]\���іマ�8Gh��oY�J�ݪߛ��Ut~c� ���������8�i1��+��CJy���dZ}���4����G��Lq,'yAE� ������N_�=w�il�4�Hڒ���W�4��3������D���\����k�>��HM	ůy����3&y����V�����S2�~j�R�?���/Q4�a�^Ix��p� � Mԣ>u�	rN� �G �z}�r��������o�f��\]�Ep���_*d�E#GꁿkT�Mq���?�a9�`��3�D��I�F;�<�3i��T��>�
<	�s(W�"�P���&�ވA�Cs�ܵ�>�>ٯ�)� ���r�\��m���"<���J�0p�L�-��7*&s�@a����m�&s��Kk�E7��Z�8�|G�zJ���u<��ϛ�H��1f
��mU��˄��~+:0����� �3{N}�R��p�U��0���[B��� �F�^U|�i�,�;�#Qo��y�L;�TV�ݚ�Tţ�������C�B��$l!�@�\��_�rc�5����@ȏ��[���f�b��M��c�������/���r�I_w�����X �u.�2��n>���^)��7������%7$9����
��tO�-�
�C��ոM,\��9�`�>S����M�$Pᔵi/Ô@t��#�'Ym�o�u,Qo>g��Dư[�bB��r���(m��ƴ�̭�}��*a�mA�>x���P2���͖1�g�G���qpB�C�����ֶ�g�x�@폛���>cޅ*+��Ȝ�7��h_�CVf�j�Qüq�Ĉ􆒐�u���&̱sǪ�H'�|q؂%|�f-(�^��m�p�R<�3�´�B}5������u�-�ш����e^�_�6�Џ��	T�i�(�_��X���;�󃕘�=�|����S�!LOs����,� �Gw9�[��L ��s�J(���{m��s���F`ځc�4�I�����_
I��"�.��ڇ�k>WF/)#�fE�Ӛ;�l����` t&=�t�d5�,��q��lP�^ɮĴq��*B�ڧ��_��9��T2�k����d����|��"��Q��j�x����6ݟ�#֞�0�M� �D/z��m�d�߶�ǰ)���� ����9(3k1`Nx�w�m=�{\d�� ��4��OU|�J�ͳk�0��fBXJe&�?���LL0*�}�d]��Czō^r5L��>⒉�\�k������3�<�͸�������/0�~�V=����BE�@=���1�:A� ݾ��g���ޓ��<@�=e�
���AQԿ����^���wi�KE��)?c�A�V�+�|��,�y9^t]��>j���p������O���$�ӤW���td> �]&��,nj"��SHe�i��ޟ���9�<��q�����.��� �_���K���Јp�yt>b�����0�1�$f�O<�6�b?���������CE���Dv�1O9��<A�C<� d�J�s��:o�f�zI�B��NF�)r��XuF�jrM����t��n$W�1�T�Yo�?ڗ-�:����?�Bۇ��?.��BB��)����A�PSa�i�M 
�vS�b~9<֝]Gmj��]��!�:��M�~�H^��Nӌ� Jz�l���P�r����&Q�����#&4�-5g��B�m\�y�{��`b5f�h�/[ �a��@�oʹD*��u ��%�.��Ϥ�.K�2]ͤ�ڑ��9E0]����d�\HJ�$�V���6�d7��lޣ_<d-�`�|�������a�8b��j���s%W�x����:U��c��>���� ��k��ؔ�Xq6��z4�4D��;2ib�f�v��/�����6�HĐ�%�{JO^��>B��+�4��������f|�<� h1�6�;�
��\��D�;�e��<z]��RB�'r ���Ǽ�зai�����ʣ�,T�'e��)/�[��{/7*���x�m
�d��ҿ��=�1P�p�HG�z�߷�����쀀��A��Tz,�NS~�:N�b���V���^���܂�Vb(���_v�[v����*n�}:?�c�W�7��}���3��&}���A��-!��|b3����U�G���Gr6끾(�I(��K�H�wh�����	_���P)��~��5#��)!�D]�	�9���<�B�#�1x֓f�\y���_�p��/��_��`%j���6�z�wr\A�FܷzN�7#�yb��@�#���x�O?Y'>g3�nP&�,�;�tTVM�z���Ձ*��[���MU��/���٫���u"�,L�U �Ƚ�>CK$D�*�@O_��P�6V�;+6N�h[�а�2����ŉ��/��"���2a\���}�!�J&"E�%s�'d�dB�k(ω�S�>G{�O�H+Qp9C��.`��	f��<F�(�D���3�^q�2��Q=��_��h]5�r���r  ����Iv{a ��l�_�. q�CSc�W�>�r��jp=l�<<Z{f ��271X�[������#�GxhwY��m%"�Nk[(�*��O-�=�؏�1k�~9��[��6��A�ɚ�L��MuU+���D2�(@#�;M_��D��CaA|����X�nsvkڡ���wYݹ|1̥H�i�iq�������cja�"�*�i���#Px^�Jj�1l!M�$;�M�Da
�ި��"'�%0"rBI�[���F4'&������LPL�cu� ���:n�]���>�D���4n:��ʹ�	�X~��׏Z�-�)�%2p�|o���Bo����<�+X�B�L`�{�&�L"Q�ٙs?��i1;FN�	�({Ud����k6듢��КjV}�m��-%��
��7�V����I�	+!Tov�l��ؼF>p�{�3����<���Sz���_D���$�ɞM�c��_e��쬱6��˲Rvw_�����W�`[�6�`d���CI����ܝS�p̃;Y����ɼ���i7� �t�C+��X�t��UJk�"�f�I�S��j=?PK�۷5�8N�ur��_Wҍ�!�a�>��	|V�,�d0ʅ8,�l�'�i�`�n_z� '�W��ib�Z�jp��z4j��DJ��,5J"G��āw�I1r:Sl'dD��~(]y��1OhNmq���s�f�%�zy�b��vYt*�4Gf�5gm.BS����ƽ��.]`J�H���sQ���i�ϯ��.�W��NA.��߱��4~e���H�+�%w���tg7�l��c�?y�ߩ�˪���G@����ޣ
�]ֲf���t-m�{�����2u�+F:6��u���tZ�K�I=?�h�>\{
d��r$�^��?����R<�JxE�41C:�Ce�31c�8�������{��Ԕ�ۤjBA.���Cr.��^�E}�"Ѝ8���@P��6x8���&z�����K��a��~9����df�Z=l*��~#�3�S)�����l.1��j�p�*���OB���dlf�N$)J*80�r1C��n'WZG��f��_�L���/���D�-��<�J������ �3���&G���[C�wR!
�eb����f�Go�b�7�չ+U)m���-����,�����PIX���	!�}J}����Z�tf��R�=��z�ͫ`"�s[��'����l�k��̎-�=��Vo�Ҋ��ҽ(ZӅX}�z�ܳχ�^}��
��Tl��ST1Sb*"q%X�D��<�t���sӷ$�o|9P����l`hīD~��ld\0l�I%/
�[y�Q;�nƮRD��:���JS�kO�����fɰL�Q����~���U_��c�:�Q��[��n���Cxh��t=gN�XOl O���r�~U���R�)�l��Y�h�����S��4ݓ(���T$�ʟ�b��3\P>|A����(���:s��p#s<Ot���{�ҩ�Z�����C	��3+��Fۈ�(�13��9#��̡�z%}*��\�*���.�dwp�l�����}#��D�.0�25y&��\��P�M�V��!A�^�@�[kH��]�ݡ~b�?�}@w,���T�\˷��Ut��'e�.�;��7]m.|��QWk�<JiP��l��4�t4����u�����\Yo
CP����~Oٲ5�t1���z���!�oO�TC'��큿0L�zᬜ4�w�-;����.�w�ۭH�!����xĴ7D�A"��f�@�2�Pm��|606���+�S��)�0�1kӑ�6A�>�Y(��Q�
H���|l�{Mc��8N�2��t@�e�V�t��,�P;�-vtc
����柱蜚��=�{3QZu_|�`l�|��.��tW0�@�q��EJ���|_-B��N�#L�a+9��?�U� Ы����p���� �s�"�}\g*K�����Z-��C��ֲ�6��󘧗�PY��-�!&	17����rS��L�N(e`�k���V9�l+*	�A�f��?����g�z�b��u��7�>�����75��+�����N��9fX�by7��9��g�劂�M�ėM�'��:�-��M�S�~y\����C<�Q�����F"/$p���4�)$�j�R��&��=���V����l�\?P�G�.׫��n`�N���w��lR���BC���4Ʀ��Ju���r2h���B��2��cKz��"i`_�v\�C/��%���k?-�ٟ�A!:&�P �KAA9Ы�2݉Zn�ČƬ�!q�����Q�w~rc�|�;ܿ����!����X=��s��܏\��i +�������ս�~�5�g_�]K����w@�]��I�?O��?Nv;!�߫�|�����U�/� RT�ּ	R$G�*�a�o�, bi������>yY�A<��#	I]k���r
1r�R�C��R��Ӡ@�hI"���jr�k��4�b�
�cld�n��7���Z������G$x�ãY��0���ToNo����<ι����x����8J�RT륰B���.��s �D����}���b����9�H��O��]�=�+%�����oTX�XI����0!4��r4S���A}#���;�Vj찡��>��0����@��v,WgN��%#S��#L�MJ�گzЩ]T_�yɀȂ�5�̪�p�Wz���Uǁ��_����Cj@���N{_x����;�oh<�A%���h��R�)6�f���(�t�~̹EVT�ˎ��o:-��&��!e{#}@�96��Io���/0�B��1A<̀=�'�!���OBG �=�s�@���c1�<m��9��u5׭�*"��� H���AÉn?�
J��Q��K���y^��WHC�:��b��?颺 �΀�`��p����l�[�~�Ɓ ۈ��E���/X�@4��7\�|�Ef�aG���EC��e`��}��P�c����!�3��DMl:�q�/�BL�۹H	���/����3d��1den>@��s��m��DrM��=�m6�iD	
�j7`|
�RPqM��N��j4����.��A܋��l	��Xϝ�z0:�i"�m���D$N<�
�*AvZp�
�<|��
y���D[�
{�;Icϭ���}u� !p&`�/(쉶���_l��ᇓ��G��3s���T����eJ���2ϱ6V�뮱�+q���^A���F!m�o;B<!=f�Y�ܗ�#���+s�T�"�%��Ⱥ?!�"��Ь4������u�M�)�&<�U�y��.���8Fz9��F�S#�:�7���g�}:Z�L[���f�:qs$�%H/�]���`Jnw�->4����1���.�QR8��?�b�RP�iKM4`b�֜:��^��5��Q�OR�,��^Q�����Vt�"����j9��9z�m�o�L�$Pn�U8�N�,��7������LW0���8���5m\B���d��b��,8w�g�uj=X�p�ڗ�Q������ϟ�����Z��j��Ҭ/~r"a��;��p'�쩗��_�U~:�%b_m^]�"0}���YTG��o����Z zo��J��st�׹-�@7b��m:�-�Zq�Hj܅)��GŨtE�Ԑ�����,�����?ih�2��z}�Js��?��v���Xu��a���5'�㭻3q���� *M��Q�w�a)�]5�&��ͺFUp��wx��k�wq#SR<b�+%U�`��ၝT[�h.�̵4�MxT�����x޿BI9�0ue��t�m��|�����Vmc��q�b�2u5;@�[#��i�?�Վ�Kc'�W���0����O�XV������y��L�}	�L�F7KT�-m䶞y􁌅v�ߋޖO믳�0�u�Q;��"�����/Дs��{��9}, [h���t�㖵(��u��L�?J�	]5������L����z��H��SX*�y���o�0='��S����:�>� �㝇�u���,E�Hm����YJ��/="���7WJ�47�B�����?5L1��G�ƞH��og@�ڈ�]T��^�#l�wO^��;��\;��q��o�\���J�4YG����p��\7�y9]�}�U� �-dsRq�^q�0u!Ө��n����i�GO�,��}��SD��ȸ�$����,�k8��C������^#[��q��5�����EX,���"�+�sKV�w9��N������E
˟h�r��.�QxѬ�I��X]������Z�W;�
���kL��
������u�_������	�o6�2k8��!t��MSB<�#�����d����u{>�=3��c��e�Zo���)�3�Ljξ�!������xm��]>�m�p����g��֓��LBI��b���+�3IK��2ՙ�Ʀ�,{��,i�u{�Ƞ mDUeZ�(1��G���Tџ���fC�#��)���HQ�r��AB��\gĢ�ε���r��(@�H�U���$ᢸ��/c��ΰ���$�9���ҳ'�L����\ ��e_=?��5>ȑؘ���j��\�ߔ��71iLG�
���Eݑ4����71C!XI��?���� ��Ћ��o�K�	�L�kxH(e��X咦���ۿ��@�df�o\��!H��C�n��p�My�W�SR����s�296�Hoj�~)�	<3� V��,xq�Se�d#&B*T�	���O�%k�)��g/��q��B�f-��A_�WkL�*��oD.i�s;'K)����&�h�d�w�>����w�( ��%/j����8r�����d��R^>���@�I�eC���{����[����v�.����Ey�;��Oq�qD�X{-'(S!�w���=�F#�2�|�����^���_2^�ow���d\�,��>c�Ս;g0���ɼ-�2��ب5WI��j�<�gW�J�)�˭Ʉ�e��2��n7E��́q`wEHVt��[���yВ��aBa�V&��&� 0cVD��;��D餓0�ú�V�\*� դ�٩��L���Gp���yٴ^��Y��-�Ci�3X�����}���^�5m����p-.��c݀�ҁ�;���	P�_Z�T��l�@����M�ik�,�cGvb�W����uh�����Y#efbeT�Uȋ�Ԥ�������I�����\,���BNa`�g�k����-꼜p�~?K���K���IQ�/8H�vB��W1�Am��fg�3xX����1���1>�&����mjlcD�A�{��C��B��j����n+<T�G��r�D`�s��|�c���_���/�/�d�^��~%�.�� ���_HMG��֦W'|`t��ͧ�
t�|V�i���URw�\|�R�xK[>
�8J�d��*���pH?�-�s:Z�Sժ�0�T���f_��D����4�?��܃�S>�E����e��*Ⱥ�O�i��j@jQ����Xg��0k�zZ���qޤ��]��|�P��i�����5i����u��(�r��nԍ-[D��K���&�fl����������)\�}].�!u����f��I��T�1�06�c5!����YWb�����q�u�8��B-����d(��ͷ׵�6�V�ǉ�lt�HC�u[[��Jɧt7��^�G�L5�gOwO^��c�"����(���m̀��K^��>`c1f*�S%V��|�2/F�?�\�{�	%UFFvL��jb���p۰Z�,�����o^s׽�m�}��9Vp���j��.�g�^ѿ51|n.�(�~���rö��;����J7�U���W<6W��6��|�t�6D�5H�m�?��5Ҙh�_Cr}���7��-�Yc�qy��\]p�(é}�ӻ}�Q�Ͽ�r#���OBV$o�y�߇�憮�&g�t;|�R��ʆ�!�blO�v��о��� &i*\���Fw�4����D'������!3�ɶ�X-�o��.�]i�6��}�5m��㮤�&Z��Q'��v�)�VMJ�i�)j/Y6Uw%6�%X�}ߢ�����7�/3c�U���ḯ27&�i����
�q�S�(�?�Y���&v
�|��H�.h=�tڱB�#�y��l�Nx���3��k����cl�:_���kx��/a���Ⱦ��la}_]OH(�AY�;���"�d���3�N��+V�a��#�%��5&q��c�HuE%�2kۼo�m��:�!�E������	]F�Ėh��� )ef�-���i&�4�p�Q.O��Ӆ�1�������㉾zh���٪B,�����EY��t��|���v�p)~C�LHպ,�B��WK1蜩�,��<����$�:}F.�b�g=�>�`�4q�ϓ!��M��Z"L�� <�0��{�p azFӌ̺n�	��RT|*E��S�?��
:K�m�O�0��QFp�F#X5_��
��}C�EY�����N�ZW��R��҉{�T��&��&�l?)Q��^�����hr�H�Ծ��i�v��x�%�Y�^�]�Eիp��������BK�� ��Hkˍ����&!x��=�*��OsP����	 Z�`oɦX�8"��kO��X���g���f��GY&y	��´:Iԍ������X�\���ݹ�f$4������|�j�L���1�B?��,B�)l�C��;���ˆ�|�q�-�����u���uP��O�nCSV,�;�*��q�_��[\�V����U7�K�7�ʑK�s- �d��s>��r���P�{�g���m`��Q߾�M��i�������瓖i	ߣ�����<%qԃ���_�a�S�������>fW*y:���U-��Q�&�Al�M�Lz��:�Y������b�&�e8x���O3k�`��UyW�aP��	w���e���y-�B�a?�>)��RT��<�l��ON �' ���`Գ�9���P�aě_�J}�M$!(�C�wR�5�n���vY߿����NHR'+�7�tٜ���*�����f�mmވ_�o�bF�Y֚�z�(���0Ac��=��$f���������i% M?[q��?�8����n�\��d��$�^�[W�R���Cm��Ԅڨv-�J�s
�7CƝ]0���k����^����@�uy�����V��K��ng殲&�B:�������@�����F�ˋf���uE%5�м�3le��8>��q6�YT6��I%����w�ioZ��
}���f	�g�b���;��`bݨu��,̿-����c�pB .7 � �2�~LU�=�a�v]<���k�d��������02�H:�V#מ��Ơc�$��˃Q�/]��7T���W���R�˞����S�:�j+)���/��P6`��o_i����s.��&�Ո�����WЏ}��ޠe�U.����t������1&��@��X���(�Z%�B%��M (RYJ(���z���v��*�1��V(�� &ONR�w�$���|KH����~5L�/�f�JmW?DӹN�y��p�b�.�D��h(W�D�G�x��p���)W|:	�gTO��T_�v�)��;Ͷ\B��ѥZ�U7��p��=ӛQ����۔d�h��/�QA4��5ؒB���cc���0�l�!�g4��D��<�!��D6rvr�;d�š�V���M���w���p 3���o��Kn�e�1
!ɛ<&���>�Z7>��jO�V�@��M�c��S f����RuX3�T�˯�r���ߢ%&�C޺U�tՒ���0��� ���ҏ��"��_��b-}�GxT�8Eo�D���<,$S�,`_��d������y�L�F*@k����
��"ڇ�z�=�T:����㕰����-F��QW.�"(�[�ux��]�V��鼬�Z5D���"uP�nr �H�'=��ַn3
t }dLo�2ǁl�[1Q �*V� ��Sӝw�ʧьd��\�;�E��E�^e�:gr��-,~e':(���,����/����6��m-�U	 ��
��",��zI�)V
D����c	�X���w=�Y�@����?��V��j�����3g�kǩ<\�Ԟul>n�Q�lQAn?��;�%�+��br�
���O�:���#|ZN����*B]�âW���K��mл������!���.j&vdK;M��F��9����Uv�;,�}~Ʃ�w���0U�H�N�������|�9�M�.��{���!ۅO ��@Ra��a�>�N�J��`���ÏBs��f��س����%�z��X:D#F��O��ϷQ5��1�P��wX�Q�O�y�B���3K˾9�R���a�Wku���_Xm:�ϰ��;���l^��D
���P�����i��a�=�^��4�	)�
���Y�w3��;��.�V"�sx)�e���+:�\�]$��:�f��Q��T|sג,�Yą��1������&A���A�	�G~�����A(ފ�0����ؔ�d�&P�䡂K�������?�h5��`�~bU�(�w�t��W�x��\M������r���	TANQ��i_.?E�5
�꠿d��e:��Ƕw�����I�����?��:�~��k�:��-�;W/JH�	3O���"6��=�!G_�w��`K'�ew�:a�A�9x��j�Q����+��Ǻ��I��k�7 �';̮�ő��`,��G��Cz��3��C�� �ߑϠ
�t�73�k����^�Aܠ��F�������=��9ВM�'�㒭EtEd�����w!�sq����~s��1�0��ۭ��9��.B}��h�n��nN�4G�9�3�Ҳ*h��S�f��awow*^d�<�
��Q��U��	RqX�����{�<��f��_v�P��A��矻�[�d�XhP��>�/ƾ�@o��!���:2�ܭ!�h';��r��r��a���A�w~���DG#D�=w��R�j���y����G@\[F	q��:D+�G�[��MF1䥯"2��ŢA���ֵ�O�,i�������8ۥa�-Sey
 ��Ss��o���e�I^�8���ӗu�%��A�Ǌ;���<o��^���U��+i����A�q��1eUw�1	�&�8J^x"�oD ��a�p�L_��8������Ks���"�\�%�o���\��"�Q� ӈ
8}'�	��uJ�B#�|X���|��X���H' ����֝U��pE���y\{,_�SnX7;AꢂT���@{��_ͯ�r���q�;��r8���f�k�C�(����$*\����E:2_y��.y�g� ����%W�t2���2��!�������{�^ZKB1�R+�[���P�����P��a��š�jR&9у��j(� Y��}so%[U��D�D�j^���@(�+T��jGh�0}'_+fT K�=V%���z��u��T��� ;�rit.�$�p؝îV&`5��1%����fÖ���P��r\��=u&��c������PRG�$�y�ٔ9( o�;�c�Y986�4:��p;�'�`�y+���_��I+���L���-�S�-Z�sQs,�aj4��3�y@��G>����!��{J����o_ ��	�Tu�{� ��:���Ʀ2u�2��B�G^���WB�ՓlgJu>k@��^�ߺ_�!��\&>`HtloOD��r���e�Y����~Y��6���r���i����~m���w��S��?d �$�[��lG� �P�.;�e:��|Fc���x�,π; Yw:���'⣚P���������ֶz约j�]Q�� j�}ڐq�!��	[k1�%XD���rX�o�zUH�W	p� J�-~�LZu$U���������K@�yio[e#���ev�Ӽ`�!s��)�x�(�v�%�p���v�ۙ�DE�\{쉊�&v��6�%Ur/�c��dd�%s4Nl�p �V�%�c'����p;�NӜ�60h��і@F���\�����y���`�X!]}�)����p�lB���܎V}�E�"Tےx~��Q��M<� 7o #ߠpިpZ�w���n�8�]=�'�� E�C���L��a��](`��1g�/��N!o%v�L[(ڟ��s�U �RQ�KVt�Wo� ��@:�W�YH�J�X�74�n���Hnw�[������e[*74�<�7�Z�����w�On���׻PQ�P�6��_o&�5�H���Ycs��A���_��A"�|�R)�]Ğ�<	�B�-�E����Y:d"􏎂��8�S%����3�r>,�^��g�ץ,�_k�;W�������3�I���c3x�qҚm{܃�v�����4r��s�l�|���5>�n��2�f���h�qX�p@\�=tO�ԑ:z2��uY�G(�(B�H�b&�>^ȑ{�(��5[�]�퐜�.1֤tX�Y�	o;=m�z{c��ݨue��8/��P�4�;t(Y���J��s�'!<(�{u�J5g��i���r빎������O��#8�n������13<^6�Ė}�����=m�hAR���#��p�[�Ir��G\���ߓ�	�6q���F��:b�M�#c��Z�B�����i-��(J��
)�d2��Z�6��ZC�S�!b�&���RP�*h][Ӡ�:T�'x�т��Ν��JUlt(�l�`!�����Qv��L�N�%�j�y�(��ui��S�[V�B�(��'�C$8Ұ(��G�LՂE����qB�]I0�?����|ؚ5K�`���@���괼|�5x�D�f38�eG�+�i	�D��I�O՘�ʱ2|�O��U�~�/+N����m�k�T��3���CY�F� �d%��E���ǈ�	n{|�l��VVHU������`v*9�H��Jqϸ��� �v����f�ѵHX�C�z%aIҢa��c���|C�I;�}�G5L5�2��f�q6�߮��R��!}�0�8��߽�c)2��	2fXEpR��:��l����Vr�띸��IE?1�H��6��h�T��j:��T���U��O��5~l[�|�&�k��(cŚ�`ѽ�a�I������HCe���;f0b<�$��Ӡ.���8�:�R�أ�%��Ey��!�wY��
������m�B�aX�a���B����{R-��HwR�G.����c��nL1�bs�^+3L��v��I^�E����?`�v:��#�΅��O/B���z���8st��0�G]t/�c=/���֐f�`�hl�*�ɡ�ޞ�@�3cr�N����ڃ� n��X+������led�K6m��u罌~ʉ�	@4YS���/R�.�T��Yt��5=���A��}X�C�uRl��5�� Hg�
�L`� t�vn�6 ��g�O�xŬ���W�u�����1af��yw�K䘕���D�@-��&F������_���YF0��~�ݓg٠�o�dT�4�U�#G�qɊ:&.�n[T#��N��`��4��I�i��¡�X�!������/��8Y��%q�d�5�V���>�
�W�� L�b��C���o�B�W�v8�\����e��T	��K=O����LTwΫC��;G �� ��?˪���\dJ��Α���3����M�m5�M8�i��"�݃w-.�:�\z�f�v���F*1,cP�!`�{��\*�R��`�R���N[F�����&���Y���n?����y/���+����$i��Φ�pZ���ͤ�7��b���k�#���}���ǣ��I��/N�d�&㥬�:�H&[Bs���?��5bŜ�[wo��&G���T�v$�Km|�%�w}|^�u�x�Ń?��P:�d�PN�i������;:`zKB�����%�6���`P-�3���#��6����w?�� �w�:&������5_h�F���N���̇�ЛA�#-t��7,�P7���\X��[,I,�G��X���[�t\�������"#��\�����D�OT�HR�O�p�^�0��#������>Mz�ǃ������fm~�>z���g߻�&��E�qD�yK@K��� �k��2���P�寡"z���Q�u�\���v�ubX E���G(�����y�C��K��8���%��z�}����͛ �	;�̐b7�� !�$=��������gz�������1�l0V'OD�r�.��$�����({ϘaMnZ�#;���n���T\P�!�̳(�"崩�D⹔
�K-�	�ݥ�y�A7!@�+�����.��%�����%%*���e�?T$W�����K�M,�7X��L�Tۖ�Q׉��琰]ߗ����P}a���M}���*S,x9�?'$e�^@58r�f�����ꒈ�h^�>�;���< ����&�ÚO��nhJ���d�M����,�D˨xբ^`��bӇ<¼C��?��D֨��M�9��M���K���Zz�A�ѳt��)}"�\�b�7�cW*5���?�j�'9c�/vl�
i��ڙ��.ξ���Vb)������������1���+;�W�E��	q^o�k����Ey����ɋ���:Β1k��&bX���B�0�=��p���E�* ��1Z�z�`'��G7< �>��~�&,V�蒧�K*��l�ܥ�:Ȇ�l������Zrς�H���Zob�[]̰�Ӥ�)7�zs�Dį�P6�}���h���ڙѭ��$��@أ��2���o,F55,�F/�
8��V�sdUοM��s���)����19v�6�F�n�� ���/R���CJ+���3L�N����g�m�i(�Vy>�����k��H	�S�`k��Ї.m�{dt�Z5��ͱ���p�K�'�*e�j�.�~��U��A����-mw�s�4�%���i�\���Sh5o,/ɤ����x�^�����cx�Dy�@H����
��撍�{1��ڋ��T�����	s��l�A;��Ѵ"sCqH��mЭ,r�Hw��(��e�.�2�N� �WF�ya²M�1?�hZ���� ��w����5��T.(>.�F@N\֯�ݫ���dʐ-���]n�_��!�g֣��R�O��ɩf�$A�S�#����Q3k�A/��T}ȑ	>��i�:/6�c�>�g��%g@o�d������6�oT�8]�BS)���O��[C�E��w�WVJ����o�L�Ќ,�v�;����җ��b�"%�A)i�9RBI�<P��)�%ܘ�X��ȵ�L	��{�\��N���h0`C�!��a�����O��B��>0�3Ԣ�bP,.��$�pw�^�k})�#;�',[d��!}K�{
�&HA��S+p���a�Q�o��!��ü���'�v榸B�[�q<8m+J�$��r�`��d�O��~ۑ��V?A2q�h�Q8���tBye�&+�4�%5ӱ�z�ʳg�F�.
{#��8J��^=�������m�5��Xi������B��ҽ��Mw�~W"��`"A�O�?
z�O�=d���.�Us����Sj&�|��"VO�Ӽد�9�k;*ČD�3��2ȱ4���E��T����.�"��_���g���x�3�6=&����~o;V�J�������8����L�d����=��[��K�#f��3��� ��]�d9��e�+O��}u�6�/ߴ!-���z�)㮸J�O��US�8J�����ޏ���ڒ�:5h�U�u��hc�=���Cj�	B��ӗ=��/FTS=��h�8���~Y���3Zhq<�Hg\��x��kP��s�s��7{S+t	�Q,S�&e�I�.�C;��M��3m��K4�ݜR���S�����UB'Bҧ2s��v�D�,�]���gه��'BZ��W��F&��h`u�AC� �7�T��_�;]B����N�c𔒌/�y�%��ާ�M��)�AO7��*,1+q�{b��gѢ � �r�+XY=���R.�\�a2���_��YE�xH�|���Q|[�\�w��F�� �ԤV�޽t+�pqW�f���<J��e^w�X>;�������|f`Zfh�Y~\�v�I�-� �:��V��&ܯ�$ŕ%�K��|��͉ց�`Q`�/�����Q��@�V�%�IJH��:Is��~��i=C����L�R�z�G��=D��r�񮙫��M��)N����)� ���[\��;�t71�w�!bYl�O-�[z"jq�+Q��km�Ƭ_���)!|�����*��1P�_�e�b�r��?��"9,���}sXtW��B�R̯�`����S�� �Gm��I������ahk��{���ZvO���Ǩ5�2�5���犧�ɼM���Ҿ�/�Q��z�h����*�+��m��jr�+*`M��v|�јL�q��v|�.(DXw�h�"~MPvG�����o����?�&��Z�rl�jyT ��/.���c��-���+���!r�`r���O*�{�[�/}�}��T�y�c���*/�/�f��gY��x�d>��.��i�k�(�!�������VS?�\i�f�����?���OwI�4��ߵ�1���F��NMT���O:e/{�B0����SN�ÿw��@G:�J@T�{��"�[�}s��\�s��j��RO2�~a�_	m�3�s���g�3�YP�n�]ׁ����Aӽ��2�~�#����,[v��06$�"�Q�����܋�����*p�qX���r'�=8�ב)vc�>�!�8=�����oE��͒x3v��WpR�k I��'>�p������yHM�pD�Ƥ���az����;�|>#�ԭ�DO��lA$w߭�Me)�Y��:�h��R�1p!��2��ǉ�+)�;ĉRQq,*V6�Ng��5�'�Sl����N���ݴь� ��n�dg�C��� ���Y�YM�2�v����u�o��.���p�~���+o��I��k���{�|�|�n��vPT��r��,7I'�p]L�wF�A�m�<I�C�rj��+�A�C�	���]�(�
��ζ�u5��P0C�J�k�pZ)���.��U9 k��V#pݏʖLՆr_6�uG1�kc�H�u\��&`[�nvѬh!U=�Z�T��5A��8g���R�r@&���{�����w@w1��� fz�d��\%9�Ú' ê����qSh��x}-����@_�z���Z�f�p�~���W'L���F�uuSܩT��V�N�ߕp�^l�j����jB׷����c�'�����iőnI�l�����G-�U�a�Rqx���A�a�ɉ	D�\�X��]�څahu8��'ɒz��O؝�>7���<uYˣ���'s�$=�كH��fB�!m�m���Y����E����I��9u
8[Fezq���I2orv���IRG,����_L����⟹뻁x��~�̼9�ª��l��R��[�{��������3���A���Z�� ��(�o�D�q�����Z�U��h�0�)W�X3}}��R��+ˍ� k7���Wǘ�zl�pS�7��JX�N�7��i��E������B�YK=�x��'r�@�-����]A�[�yn�RA	����ק��cR�/�Tw���|�؝s�����(Q��o�\{���.��F�#���aFsr�X�S����q�.�4;���ۓ���<N�o��U�����H�8�W�Pىևqb��e:���ۖȃ����s	6#�݁L���FُR�����q`��[*�A�����fy�
���T�C5�q�+�RW?1;7,��c��)�V�vU��&c��9�"M�iWEWJ��¯�yV|[�嵤�<\h�E��?@��azY��S�x�-�v�:�6;jQ��2O�Ď���?�����ϯ8�d��I�$$E������A9u�g�-J��f˕�y���4s��%�z$^�y�����C�Ac�buYt���X҇�S���k�u�L��׌�Ҫ �/�h�1�ʉMPK�@b�$d�C;�zQB�(2��},�J؋�',1m�C^_'=os�����sP��?�4�DP[:@cm>����O���;��7���N�iUojn�',.��o���L7)�lL�Z��~�2��x�3.��Rb����	�#��<l���p�4}v��J�"��)'(�2��I�7�_U���f3�;��?��5��N^���_�e�h���;��l�!��1��H�%첼7;e+��W�a��qX���A����*����z��򡙈8����]I%�}^�R���8���&�eC�;��C�I�-������ ����<�G�5$w�Υ㕂���*�6ê�P4F�p3���_k��l ��"v�v�|�l�r뽸��՘f�%�Z����W}�<C�?i�c���e���*���2ǅ�nV��`�Q���ke�\��\�w<��!{0���n	U|������Z��V3�����.�Z�Ļ�礻�a���+K Lo^Zgj�n3�#�[ *Y����b��f��lI�D5��#�Wi���$�t�Mc׺��)&SW� �p~,r#{z�©�A_�zIܚ=@�8��wy�����O}�DJ��"a����T\���.zN�~��	=K�YY������w�ָ�s�/��������G���Pa���¹�N���Ƴ���l��^M��F�GVۀC�Wtⶫ<迢P���u��o����33�[`����`o:ǒ��~ C�O`������]���W�OТ��7~\�̾��0����_�+f�z��=8�!���2ĳ�u���;�ti	bD��ݭ���+`�1�"�(K���%�;1�6%�<*2'�?V��;�E{��FA`��ʀ�`�VӽCÌ�=���q���0���_�X�����wg'�q��qm0�KV,��촖�(��� e�%��&��Kov�����*,Ê�!�$�;���s����zӜ�.*>x����>�̈D�T�V#��r!�?Q_079�2�ϊ�����xfn�ܒt�9���H]�:���3�eg+X#��͌(̍��x�R<`��
}���`F�洉{�a?b�<R�����I�p���W��SZ<h�9���Ƨl:��mt�3�!{C��0Q��~;���:Rh&gAvI
��d׻U�0��5��_M�<i+���q�~���٬�&76�p��o���d�@�5�����f�Հ!�xH���~��!�P۞�4�7�@��f��:Θ��5Q��R$��\ɑ�}h�v	����z�W���'��%H4^��Va��1ݽ�y#��(ɻ|�ӛB�ZB�Oj항
��.�!9T���e������,W��Y$�Ⱦ���^\�H�@�έ����L�g�w[{�v�p"�q�x�pe��������!L���x��/2���'�J��V�+���,��V��!\�i�{���[��
��B�	�Iͬ��n�������b��d��[\���O����ne2�L`�d�#��R�Lܢ�hˡ()��j�� mN�3l+�@ ����;*j�D!�W�20!)g��S��"�H}-����V�-�6.�����BF��jp��K����O��g�.�#�l��zyfJp���ޟ�W�����˭�C����uw�&:�vދ�՛�%x��������L)��;�;ۡV�y��G,v��Vg{�S��K���ej�u�m���2��_X��]�$sw���_�m��:�T5�R�Lg�E�_t�g��!�a�/�������%�O��*P?�9��÷TJU��ՔY�E^ID�^Pa��N�����M'���@�e��-&�m��/}���NT�,w�tq�E�ڶ=�GŜ+9+H`kG�jVi��u�N������ViY�%Y2n�w�Qh|�:g��D��_E�>�����8�0;Ma8��g��p<I�� ��� �����J0�Vh�cJt���S����Z�˂8`�V�A$��cp;J��-�حF���b|.n����Dx��-&��.��Y����қ{�-��F����0R��k�srM"�2q"��5�P�a�,�%�6��N�_�1p9���r���q!���{h\��s���$�//*N�a�����e�;�v��C^�9~�\<��f�l{u�sH:J[�x�9yY(,xˎ<��A=n��}'��3�St�t�Qi{�Œ^�0�C���+ڐb"���DWZ�Ľ�Y\A딝@�?A��]�'�:�����/��MjܸCCo��{!]��Tg�X3�i�ܽ���A�a���&i�}����>���ho�|��d]�Jq�<v�5$Hĳ�u�&�&y�F-�:37J���C�͂��̅�?�H�1Ф�����LG��~�1I{֟�z|�J?���v��o�"�.�MjП�L^;p͉��y[��aȑ/��pѲ�?�-�p	��-��jeF����J
��۠�O��w+r�&"
R����9�-���#��<�E�x��@�b7��73ILWjN�:����{E�rʽ�DƼv �� �H_xTq����	�S���.�6UT:7k=l,�%:��!�t����XҤI���^�T��;/+�A���{)˻����=�Xi��Y�j'w\�������? QR�8(ߴ.�L!;V��]�@8�B�(�S�^о������4Nq�\���������C5�Bbgt�OY5U��_��%�b�*��]�z
�����x���15�c��=Ԑ���v���j�TW��ߣ���h���/"!�gpDWZ��g�
3��|��VH���sP����M�mu��������q�B��Dd���;�(,,m��YxkӘχ3���d�q�Jԃ*��_9�U�'@\
8�fޱ�$3�����-_R��kr�,t�~�����oHÅ�	~��Z����tr�m0K�d�?]�ob�*�U�GuW�Ng5.�;�;H�Ƙ��F����	%U��﹠iս�*�OvqĨ΋.Bn0�}�K����a��÷��$ִx#U�6�؍�o��l�3!�~��`���G&����փ��?{5�d����}&���6.coRO��U�Zby@0H�}t	��Y���{�3=��7�
̅T��Sϣ���܋�����"{�f�T�]c|I��1�l�w���dP�/�#�%qA��Y����4�&�!B�c��OMԝr[x��?�S���+�MJ�܆�}[U��Khv:ѡ<���^�2 G�㤸Fb|*rR�J*=Z��ޯ���ӵKΪ�8�o�O���8�|���I�r���"�}�X�6���Wr]��n�d�a�Q�� ��Nw���޾`25�m��/�:��m)
2��"	 ፸��%`S�0k�~O��!�v��	�pM�� �!���i�6c�%�݉��*?ak0�}P�����O�JZ�x%/�����x����R�Sinv�u�e	�5��N��h�\��ݑ3Z0��~�jaQ�
W���8���9�F�OH�t�
��j�/X�豭��c�;���вIt���"��	��ڈ�����<WYt����8�� �'3Z`x ����AA�	�!#�}G��}&����#{[�+%j�7t��Z�*��'"�z88w9"i+�_��Ӈ^?����y2D�	�[�B�ϸ`���n��kOCC)>Z������&0�j���t����J${Lwŧ��������Y�H1>�Z�{=� ���h�xRy��O ��S�h:|�<�����{�R�� 7(�+ۜ䗕���/��G��ϵ�D�[�|�2���]P+��	O�Va����;�M��/�ar��U��Z:r�5��i��IAl�P���и��3��ۢf^����k~�����t��O4���<��Hpݞ�=��)�y3w��
nMa(܆���G��a��\%�������I΁吸���c.0G���0Aɿ��/�U���ʀ0@�+4u����Q�;8M��Z�`����D���`�O�Oe�(�Bmyd%̠���<�ȱ�j5�A��c�Hv&��L��w�ҝ�n�Iv��7O�mEC��Wd����[�������
��O�0�,l�f3�t�j���qG�����W�Jر�|n�|�~+2�#�� �	���gQw��v�v���sP;���O��c@�c(����������bf�b�C.b��&�S^��d)�6.���d��x�epG�B�'\S*���;���`�,b�=��fy�nW�oDa�.��#���s��)),L�7`�4�C�^3�n�Z���Ϯ�L �ҩv�ʌ;b��:����/õe���Ok����j ;P�|\*�nf���q��m�%���^�K�J�K���#YUl�܆�@їh�Z�kA*�cd}{�9���E��Ħ�8\��M�o�-�Gd�N	�G&hJpo�pV%�����&��ds�İ��jw�թ0�=i�Jb���` us��K7�8���)��Xk=]ɺ�faw�$��hB�w��G�#4EIz�J&ϩ��׻d��S��A�h��X���^v��H �&���Ͳ��)��pb�Ru�Ǽ��¾B��Ez i�Dji˕�/��0��8��_����#� ����M���!���� ��8x$}G|x5'��w��U�����Dd�R��1bkI�{y�*���D�M���`ݗ<<�7
��˫���zJ�Oz�;�¡پ ���Č�7e����4OL�����/�3�`��AH0�����#�m����*b3n�fƁ
'�!oJF������t��������3.��Q�܏^쟈GyT$�f�E��>>
�i\�e�CB+Bϱ�a����'�Δ"����sPI!*��=�@[�O|�@�v�D8��ԡ #[���d�!�2�z�­E�'n�]p�˜�7�p�u�:ikӇ����\ȵ�k��m��*9�
��;�� �-���0��HokqI��˧$�=� ��Lt�f�dl>c���?Q��G�Q�P%��2�,;5̫��[$��E��qP�n)���Z�W�w�g�vu.�h�F�%�Y�:�JpJ��ʘ�(�êPߝ� Y�}d��s�>����o�Yz�Y~�W����O<���˪Ua�
}G����l���${TP���",ds����֛f��i�+rBO�]�g~�^�ֱa���a��;J<�gW�
����#lk|\��,�aIO�6C�p��wf����d�L��p�OsK۷��\�gG���aB�n�+5�E��D�M�����APk �艕M�lC���J{�%����o�T�<��sR^��~a�t����Ԯ3&_�/*�J��DK��D�
��B�/I#M��6I����i���,����|����C��H�zЃ=��]x�����ؐDA��[|�b�����s޿�t�=������?m��걈��@�������|�$=�ܖ�R6B	h�A�4QH�lUKJ\:&��y���Il����υ��2D�� ����R�RK��.���:�$I9[��
�!v(�H �,x.��o����^��~5o�ꂷɎ�ʛӄ.����`���9'��D�×�¦�3<��w�O����@M�^9��V��/��"�nSfB�#���=my .6F�
Z��<��ǳLP�.	f�Ⴏ ���⏨��[:@Tz.�7Ú�C��
���e�s#< �{ťb�&i:�+F̌����%L��<�8S΁�8��?�5NG�H�0PC�W�H��������к�����a@P7�C7���3�^Kq�FV�|号���͍�ƏY���HZ7�	&(��1���,5���b�xm����b��@�΁U U�Ei_Ǚ����]�y$m�dO ��2� �n���a(���+����r���,W��&7�z�7d��١��~2�11���5�!M�rLE'����7�,(�կў
6�Hs� �^"��P�'��E�'�?��
RB��.p�`n7��Y��(�i�I���� ��u#�y5b�_,��Zb �.�������.<�)�� �����i>��U7��w!���ꔲ��4�l�������	u��=N�c�ؙ&a9�q1+����+P^ް=����a���4c�&�����ʘ�׌��׉�$O�.:�m�$��q\Re��W&7=DE��%���kny$�R;�OݙOçUdL�}�͆�<���@lA�`0�	8�勐�W�J1I�]g�G��'4���;�����or�(=-6��W
�K�S�J�}��N�|�	{^$i\k���GБ�'�;��kg"��h���K�q��%�pf��vP�F,��i��w��ׄ�͠�dױZc�$.`��Xq*!�gM{�:p��B��G�݆C�E%1X&��o�/�dOL#?�i]C[�
�+*-�W��$��_FP6���ˋ��d�L5	�L��_�0O�ٙ�w�·a���%r�O��4�` �⣄��Bҡa�
�_<PpL��L���Q��Ý�E�1�K����3�=����eZ��7W�������C'���� �+LU]�T,�����"���!�-�GP�.�Fڰ������B��`�d%5��b;e��}������A��ɛ|%�Gs拦�S"xR(�A�C�OL���!����2��U�E��w�	&�:����d�!G90��u
4Y2��TI=��Z+����FK)��������3e��J�UD�����8�;��ӳ�_{�R�wUA�T�lJ|�H�O��8���rK�w�^�>z,ވd�/�Re�(����� Z�s��wLi�7�X|84U-J����ᗼ�7=��;���&���׺�*��H�V��`�Fb'�dR�(0�Nj����9!�?��!���}ň9;4�Z)�ּ!�4!m���]K�Ĭ<�٣�V샤���Y��fzi�b��g�i����j�0ꑝ�H��ʙ�6g[5� ג*ܦ��G>���eW���X��}A����Z\w�X�=��٬
���I���l.;8�M��?�V��n,���<ՠ:�H4�"���`��O���Oʚ��4y�P|MǷ�95+Ilfľ�A�a�ƅ�+�50^�'�x��A�X�$.�''`&��Z�g?e؟�J1�d�!ydϨ;��N�`��e�y��Ꭲ,qa�N<�>�����y�*��� ����ŝz���H��1���Μ|��HLqxp���n��r�y��K���{����R��s� <BP� �"�U>�bGe����:c���CL��K���C�d��V����gH��I�����;-��"m�p]�`����H���)ubN�w��A�o�1C0�;gș{'�Zd-м��J��wG�(]�;M�ç9�]X�.����Nq4��@��M�j)Zڳ���=i؀�A�J��v�5p����e1=j6�f�쾦a0���-2�l���;U�Ɂ�X���x�*JD�(\�Eؖ�I���ď��6�CuP�]u��S�� n#,�k$��4Yxd;�Nq*�U�)t��A�,�zv��f��{���4�{#�K��Tw�������k�/�Jv|�[�q$���!�$_5u\�R�N������L3��+�f,j� ��i� ݂�t$��
g.Gt��(QJl
Eo�d�n��q��.O�#�$�_�ӫ�p(/u�^sse� /�S熏]�[�+9g@�	حܱ�ܦ�c+�#�#ԛ:��`�Ǭ}d*{	z\�*ž J����c[�l/h5=�Ҵ���<`2���@��a"2_��D£��h���m.FI:��=f"���n��\R��Hb?�)�m�A���H:y�[ח2���/����1X�o��8�#�Hfq��_���^��\c_�J I8J|�6�����K��->�J��{@�&̇����襀e+�8�~���}��yA�>,�>Z�:��L��ʨ���6'P�"�e���Zہ�]jH�Y�����|$�o����IBu��z]`�й6��I�l���Q7�H8�{O �9%�v�q��e��u�932zqę���/��T��.�4�iC�P�Kڀa?��R�*^��{r-�|�s�|B�n����?Ca��?o����V(�uρ�o����>�I�����m_'���1��Pת�����/"��lX#��M�y�э,���mr+���E~R�B�c�E��`ţ:�gw2��
�1���Q����_�'�r��(���> �$h�f�e�N��2�NFY��Ӛ��{P{��P$)�.�>���8�YkD���0�e1<���@zZf��J|� 婁�.�SlH���զ(E5Y4�~l�ê���O5�� ���ԶI����k�m&a���F��$kל�8�KE�q���ku�i���V�ės����]���վ���ى��fG�kFhd�|) #��V�2�?��Yz�����w��(���PY�w����!���Fa���S�����.zr���]��ҹ�uL��u��o���9!�
@ܿk4>1�qp��E�%bw�ط0j7��A�=����s�����ς�J0�
a�:z�uu�F�;_ 9 #�A�t#)c��X�|���Bs�D���o
��T���%H��x$AA
1�b���oW�GIx7*[�d�� 5��L�H�H��'�İ��Q��MQ2��rq9��ɯI�2�7nsK~ӧ3��������������>i$8�,�|�T1�e^[C�
wxQ�Ͽ�������-�c�9��:�7��F1�O�I�$��$��
~m�9i�����|�ݢ�V��4}|)�T�s��2�*��N�&d���G���i�-��)�K�5���9���U͂ ���_~f%M\�ַ-�����."��� d�2�<5��Z�%�c��n�.�y 5z�?��9hs%��_|>��wJ�h���3`��_曀�Z�$�
������$a�դJ��6�d�1{�^���ղT ���`^�B�WH'����W���%DA���9�u�, i���{=� �+7�A�TVB�L��I����M�����GZHa'M�9����*V|�yl�4��	����-X
��Hs�pc��k2��;�aO�2T��(A5T{���$1Ң��.��\t�\Jg�`�8�ۤ�}?W��e�`�"r�ȏ�>�h����W���_�GM�'S�li��v��^m�q�`c�OC�f.�Ԋ�^���
�(/f7���KdY�먗��k_zq*��I���+aR��Y߃�9ȑ������>��J��̭P�GEP�`
Q�U�7o(u����e��u�&��@�Nj����NЇ6m��2���C[@���J�$Ӯ�zh�|\G���I{e�j�7����s:+�M�ߐ&���N�a��o.��5 찖�X$غXz�=S�n{@�7���Kh�ʹ��Y�-�.���hdtrۗ�$���]�F.Q*҂�OO�����ƃۆ�O�Ub.����oL�����LDe��	;�>2��L$�  �_�6�Ѵ����1g8��7��(�C2R�?�����s%LOB�������87�����j��M>��\:Zو��f>�t͝�rP��~���C6W���qf,��i��M8I��W��ۉ#ħ�*u�:��h��_�'�.aK���]�Ԓ�c=a+�n�Ab�Y ϑl�ш�0ܕ�v���֥y��WA��<���n�W�X�*e7���p^;]W��Eȯu���d�i�Rt�]7��s�VM�ߪJm6�|I_Z�/��3�����I��|bE�486"Z��
�^n�4�'�%|��̎H�D��(~$������A�F�\&8>܎��AMx�M�1	�y���)�bp��e腨�ɵt��a*�$�'�jv��������v����B�d�e��J3��	m����X=]�b�s�~v�B�9W"x0���J��d�Qb�9�gѐ[Q������E��Ъ�
v8�BS��8kLf���<I�O?����1���3����Q�c�KB*��ߴ��&q=��B�b��4߆��5O��N�I�[�Ul=ݔ���l܍�����B�\�ϕ��\�"?խ<Ƶ"Ė����v�V�|$UC]������J)O���e.]�r�i�jQ�PZ���� ǃ�[uάa����F�^�Mmr.�K{ 	��UƆr�: �O�d��:E�>�YO�����1�w�nI��[��bG	ޫƉ�yn�;(
��W��B���qK�p��Gؼ^D�^�.�vL��:`�Ҿ���ߟ
C�wK*~e^HM���!8��^1yV獖�����ϯ|J�X4�����$	i�0J��6K91�Y���PSK�5��ݢ��,�7W~%�� B�z�ł;S��6�F_#[%���7ov�_KpE�����	(n.?ö�ՂyN�3�AS�)�vi�cNgM�B.�d�X��	�D��Q�c\zO����uk5.Oj$P�s�-�5}�An3\�څ���/�%�+3��$����>Hݱ���+Rs����=J�E���l�a��.fN1���C�}B�L�ƿ��e��i/&��]�XX3ʣ>|]J��z����wG���C�姕�3 Qx�w`�o�e�s!����	�mT�e�^\�L���G}��͞�nhx��rN�i\B�a��P��0a�L��W�h`��`�e�vs�������>��Qe�.a�j¬J�zs}�m"1��>E2�{��8,a�*�k�#q �i���W}lԲ�z�"Z���j�>t-$��1��2@��Vd���߹4�v�����6����-A��m��m�s�N.��v� 10���8x�\�����`�s�/^Dk�qD�����ǟ����#*���n�(���� ��A�V׏�%i�8���$l�#��D}�T���EA�e	W�G��g������t�E�4yu��J��'���E�Lt'\3����.�LL���l1crMT����l����ڹ�I�#��,dEd�I3�����Q$]V��mK0[l��Wx�,����)����3Et��[��7k�k`�h/���H�Nߧ����sDc�N`�s��ԕձ# ^k�w�8)^)r2�.��ˮ7I$��2�#�fa��t��`	;{�d$7��Yq���sq#��d�b~���iG$ݒp�C^[t�z����̙kLW�.B�Pq]-fwz����N6�[�����Bvly�ק��[� �"!eqrGӻ�݊m�y�x9����7G�0x��>&����;�G	�~�q>`df�?ʹRUb��D�6.�û�M+�/O���y ��kv��/H�:a�"�#��7��fk��b� � r`�e���d��iӃ{ʌ!Eޫϡl"˛�Z��_g�rt�#�*G8�с1k��0�H��ه�u��;�/��s��#�E-�W4�����eV��yz<�9:gUZ:���![�a���ӕ��I�IMv���3yם�-�K��-���^�����Ҕ]�f��Hr���$��v$ֺ����!��u#�^g�v�N�9�4{����n�U��U�l0��̘@��Z¦Q��R����f��Kd.�+��T��U�S���E:�T��P4��w�YV�P(n���.�@�H>A��Ku�8�S��w��I�C�3�Bg�@�:��l�Wz��,�3
���}.�i9F4��&V�o�@s��{�'cUwo�_���+)�H(�c[96�1m�
����7� r�|zp�;�x�y��Y���3W����k�:�7��m�?��o�Ĝ���d�x���iC�S��Ϩ���	S�1�����F�s =������W�uW{��T�I���g�*������{\��d���s�i� �H�D��'�����rp�T��AWM�-[ũ�~�qSfK_y��%x�꠹r���W%@���R{�R-�*-�!��T��AW�\^.�0�<.�#Y랯Tn�{��;ӷEp?h?Ǎ5�_��/�*�)�ú�fc�d�ןnu.���=��LY��o2�FTT΍��aB������)�E�{+�?O):�}�+�|�Ͼ�ô���2h�¢�h0�T��%�4?�6��/�-`&����~v?z ŝՏC �%�%\�+Y�~�!����Me�j���!�R�ΤQEFM���mE�����aZ�K��f�1���O��0Q�U=[����ӡNi���MO.�%���)��=���x�!˽¿z��,�n�3�u�Oi��]�V��P��a�n�͎pN�M�y\�XD����%;���+�{E�z]X�;�+���p�]'k1'��b_$�7Uq�[�ۈo�_t�N�*�f���?W���w�Z�?�k�R.��m���f��e�X�T��5�KS�_7���u����l�s<��a�#��Lt���/�z�揄�썳zN;�R�!D���9�[�/]h�T	��U�z �����K�℃1�3��R	ܱE��� ��<c!�oj����S�̎t>%�9Hj\�-�^jI���p\���O�c���lp5���z��ڞ�h�e~�O^�/wiC?��9W�ԻNL��	 ��>���ǐS�/�Y�G����=ݼ4�>.>��P���+��:���A�W�)r��@	: ��!�6�J�������~c�v�|�~ִ}ۋӻ����E
�l㈆�%])���xXy9|儥d!��P��yu`M�PX�O�4�Rԧ��*�����e�y������[��"���fV��6����6xL��-��tj�/EXq��|R�ژם�J�>���*�g�0;��Pz~zO�"�o�S��2"0v��!.�p�s��9PL����Ա:鏃��9녉��Eb�3�҃�wKЇ����<�6�8:�AKKR4(���[�A��@K	���ȳ7����L��YA7Yc�Ԛ,���7^��E�  Kd�����I9�4ĕ"�Uc������e�$����H���Z�VɎ(�Ȟ/�Ӿ����ș_�EU'�<�c��ugH��\�p�����$Jv����{�'!��S�䭳�56�{e}C?���f��OcΜ���������-Cv��Int_��\�|Ԃ�;�0��b��@l��.LW�{&����C�$a]�ٟO�)���|�p�����50��K����o$qGv�%�l쎔��=��(���/�ñ��ZV�f��1�k�q+� N�_��p�a��+�p:
c���)8��֫�\�^ܐ߬@�b����X�hk}43!���o�wyF�1���%t�$lmS�5\~	l��6T���[,�ݕ�kg�3�C��7�g��D�w�R��g�e�����>r���ͱ�ڗ�q7�Mɺ���0�r�\��]�=/�G�ou=Pw�������3Î��i��)����R_:.,_f����31!�R7y�U�~^8�5�dp�����)��t��k� gp��#WYG��)~��|��H�u�=�%-!{�)�;�",���-�3u�zPD����G��O5�~#��#�/�©(M��t� ���)J
�R)/�������%��� ����P��.$Z#6��o�����2�1:;�E +�#7$���K���}�[�=,�b�u�ӑ���`x��'�s�(Ȫ�k;�p<0>6������=���2u�����q������L�A5��G����6��r����^z����:�c�(�sP>�w�G!��=�l�+�\���`9����B�CL2�g4�R5}k͙i�hF�� 0|�~���y�(g?�/�+?p���_��Be���|m�jCI�:j�������nⶠ:����!m���������E�bť`��p�w�pd�LE���*\�Vy"3�3A�L,(a6ȉ��x���"���r2�P8j�2,�q<"OMP��d����p�g�j����$
KfA���+/bM�!�Ut$�N�l&�E����g��^�B�.��sZ�V�lT���/~���?��$7̈N���z��|�R�Rb�x�M��{��N�B�\�9�T��y��\A19�=HA��F�1r ���8dHn� �@�/����+��"��P�1��� �#�lĹ�Z�������e��ܜB���=�6�#���
��&ִ
���r'�{M|k�VpA��K�++�B	?z,��2_�c�����l�=r���!v
G�O@΅�}�K�"Ӱ�b�����д=��s6���5�x#/���_$|ծ������d�Ex;�}NBy����c�mVe}�~��s�}�͸�J�wl7�W?C#��R�Yu�z���k�n^є:��N3��"������n��+j@		Oo�OS�Zq8!��T��m,��C�F�,:��5a�#S&k����1��x�d.��S!�2GG�!�{ Ӳ4���#���n>o?J��x�	�Bp�
ؖh�1�'��M��!� f����z��'�&K�W���L�1C�wD�Ji��DQ���Mu���l������i�!$9]Mcx���2��M���Y�{�(I��Zg��ݖ�,�g۩(�~K��f����_��ϛc���Z8�E���T5d�!��<��~�ɘ�R��+tɦa+�(Gِmd��rg
g��-�F%*�g�Tgx��Y���K��d��^=�܉-�n��D�tA���?��S�eFm\r���8Afck��E��6���g����SH*�ԙ�����2ٖ��-h?+(4w* �3N�Qw�n��Djg����	�u�ѱq�=@�Vq&�em���Z�9�$fX@�E[\c�k��'��'��x�F�dhX�#W�Դ��� �ۀ�_w����D�	�gp@���S�6m�����f
�ZPs��o��
t�E�A��z#c=Õh�0�h�j�݉Ų�i��2|�6��,���m?���Xe���[ܼw��K�h�8z*�D��(xM���ҋ�A#��������2��������[]���I}M�>�gs�-��*����ɉ�������\�S���5��r#%�w� 8!��~�a_��s0v�iRZJ���}?&U��nc)��T���4��3{w�x`�:b^������*�|�,N��&�_��1��뗚F-�qm�Z��w�D�����j?%l�(�;:k�{v~�?qW�� +0��
+�Pm�@�͡G0��
���Y�� B�O&En���t�z�W�*�$����R��
 �-�vxہAc�xق�Z�_�o��Kd�b��/Eȶ�x��'������@�#�$�u]}I[��b��N���?xk�w����!�~��^\77�}�C����h�"}t�>��0 /��X����gg��3�N����Bʎ���r�&��s�1��/k���t��W����ITq�}qλ����F����_��G�?gVQ��Z>�۠I	M��EQL"-Z��2b���X+
�"��"���(~�R��,�I���T�+k�)�\	�<����oZYW�K���Zͳ.��$�Am9Se�o��ޏ/B��8;Ԃ��l���b�\ L6�a��0��!/���,�|�S���rJ	���N�~�*8��7��������� @�0Lvf�®?k�^�WF|�[w�I��_@�^�;V��R���a�*�N]}�H+�d��G�y���CJ�W�mK�TRe�ah�{��'&�|��PGj.{����X
l���|!5���	�m��>D_��p�#��Ք�!T�Ӓ��q7��K��,�kLx�8�FS�����ұ|�$\-�K�2��('�Ζ�Y,f�WPTb��7`��g�' ����������E��O�	^��c�]l{G?N	�R7�q�"'�uqEJ0[a�2T�:2�L���y��Dr�(u���7�_�.s{�R�込V�c�i�V�9��	/2�K���
��s=�<�D�e���2�"�L�7��<q��EJ��뇨�c3�U
��2
���F|��|E�(���/E�)�ˢ� �l�A���������[݅��/��A�ٱԽ��y���y��%�z,i(R�����a�5&��bg���z�"�˼�H�)��hB����1�8@s?p�`B���� Q�� ��Gzl��T�M�:j�_��y��L�O��8̞p"�9^����=���Hh�s�{c��BM�m$�w�"��h(��-��犵�J�+.�ʧ���I}���3y^��}����M��ޤ�ptN�����O��>q�̈́斉����>ŗ�	�.&~ˣ.�kr������������Z�(l��Iv�pE�{Ͽ��#�����[�J� l��r��
Ġ�(|�q��d���<���Mo�b�4�4�x��cc�����2Kt/�[���b�0������?��i��0�0��qW�5[���Ƀ��7P(����P���Y����<��|<%��=I�[l�niD./�Y�s��+1񎧐}Iw/�>������+S�<H�~	�L-� 	��;͠ɂ�f��i\+���k��{�'"��j�{C�w��l1����oŽ�c,mh����䜦��L�߆"�?#`�D��U�i|z�x��K���O�;���㈁F� `&E{Y�.���H��`���%���}W��˗���(U�mo��g���q���T~�Lٱv�k�t0�
�]��e��j*��j�a92�Y�s��?�p
.
PJ�Җ���%��K?�G�>���� �9>��
]�E>�L��F.����k�4�(��L�?-U�Ƅ�{�#�k��I�fgn!U�)��5�Axp'Q�L�s� #`R"�lm>����I�b���00�I&��a��+cS�m�J�qZ��"ʵh}��j���CK�P�pnQ�b6�]��r-�O�6���=��4���;��ث؀��H�˲L�@�<�?,_�P/~�q�m� ���.�V��WGi�DJ0��ӮL�҆/�K��d��KM��2bFGG0���Pk?6.=�А�Ӓ<�@2��Ǝ��9d�t�2&���&�>r@�^zuZb;?��Q������l��=Ą���Ӽ�=C��ښ��D���lx7w p%�C�!A�mz�@������ݛy�P0���4�b�B�'n��-y5��.�K5�`�#�C\�:�R7�/AR\��#=G~'�>��c�G��/���9������^ø0� �hS�=_9Q;��}d�w��!��g�ƢB�����I[Ǒl�{Ai�vL:���#x"n�K��)ڽ�"@�������G����� BGWX"O�A{�����;��X�GVL���&>>�h���<"r�?2[�[>��i7I��<X��e�$�,�I��y�RQ�SW���
#�#�T�K'�wiPIDѹj��RSU�w�bގ�	�qG��3�C?���W�Y���`�+=��|L��+�S��x��7�끡�%}%�[Sϭ��7P(�{,�\4�.�AE�-u�!�0}��[u����m�}�B�ZE[߿[��Ԣ�Q��V��,9J,����j�"���ӥwn���6�_���F��r+����?ϳ<e߯�������+-Dg�In+��a:.�D;2�ū �>���S6 �^ck(_o�ӈIT
�>�9n���)�g��n���z��`�#���&{�,�lVƃ#`-��v�gR)�=7��~����(j���Y���9Ҵ9��̇�^��� J��V��yb�y�m��rK�]�������n�����Y6]�uH���]���@f9� ���q�f�e���]����N� A��uN{��z.��t�}_�7�:
:�棉`�A$m�A^��7$��\Q؋�y7�`��ݸw'8�Z/�*��Pb��l�L�CI�V�e��*b1e��w�����^��&NȧLt��%�H�FF�q������c��Mja�vي��G�3�
��*�/������騧U�v��D���'?��r|�-����[�h7�%]��{��a��x�i��6=��&j����if�U	����K�^��3.�u4�9����&�ބ��o|-�]WF�џR�tt�ەC<�Ұ��/�we���1D x]��{`���#�)���/��Y���A<V�2�J�BjM�V�vM;�NT��7`+���CT�^��.�%���%TKQ(�I��YB�8�L���Y�49o�E
9
���g~jD��Ҟv���"+3^�'�oi|Q��|����0?�7�L3���8����������6B�Z�M� ���-d��[��t���H�s��p�	�/��g��%>����GR=`�k(��~��w��$OOy3��c��Aa���%�ى�T�kh��CëM�pQ&Xc���<��Dt�R�����I?�����N��?� O[��@�RvЌX2`~�HV��`��.>� �! ��+AK+��+z��zg�<57��� ��/Q�!����i��J7�cl�����F����8�����)~�S˨�F�uS�&������ed9��j�N��ٸ����or�6��Słi:`��*B($�i��E[5vã��.��KD5)��ϳ)_�)��m��r95�)V*R|lBv�h�pHV9�PJ���#��Ւ��r�M�w�c� 5
� �S��6]�C0�R-A������/mҼ��󓚉K�I;k>��9n��H��t�K�2�'�!>ҧ�z.���}G�\����Ow���t��O)�yu�D��H.肈�Z�L3��kj��lٌ�~�]A1�������Ho�V(ܳH�?��΄k*�39+�d$��k�6S~h�@�G`@���#�`6��g�fs>��KJ"��!U�s���S�E�E���6�7�ј��iBk��ǙM1@&M<*:�f������O������v�P�5 ���2�?T'��|x'���0k�RۄF���V�/��f���O��2�.U��Q��Sb�Fg�&E��B���Lx������&�B� ��u?V��/���VSӲa���׻)���_�U/+�����
�lA�}����_|� 	^$�gy)�]��v����,/ ō��*1$g�k�.��n6����Le)Q[s�'k�<b�CnX���<%A����"���7�j�=)yq�\���T=����m����.9sE2"���7і�?�	M}��p��=c�n�0\���a��&ci%j�
�ic�6��b&,�� �wxC�{j?�զ�� ����^F-��S�cTx�Y{z\�阋S�'�Cm̍ҹ��7����m&�f���f*��:f��5��5fF��K��/�u��j�~����I�2fiثE��f�-���COIPY�˥�� y(���I)����<u��eD��7Br'`�v߫�;���潴XyŢD�6��^_"�,Y�#��'wG��`�̩��-D����4��+o��<j'(���Q�7���<晾�0'�IZ�����/����5	�����,�&f���q��<���lE���Zy��k+ˢ��Ӻ�5*IݴPu&#��i�� muyE�~D��*��fX-'������p�кw"4dݱ����.�^��!p��N&��jYx�f�,�����j;D��C�A�ް�ϴ�{Mg촕6���4>��d�}�������Ȥp ��Tj�K�987����J	�Z��Ȕ0oɶ��.�=�������&z/��}��V�!e<������?]�A�ש j�q�y����.�����{�hn˓bx	�1(s���`ʊ�"���}���ʶ�r�6��|V�H��:'�v�x�zkrp�b�X`l�"�
Č�!�Ŧ(�� ��wV%����m�cw���~��k
�N+�������~�6���4�j����!#X�qh]'�'�}!#�~��W�+���ߨӧ�����#X�^���"�Ԗx#?�bX� K7�N�`Ī���z�����u������� =��3>h��/8���P�3�;'(t{����u�<1,�?�(-ˎr���B�!��l��W�֛o�W����kw���7��JM��<v ����4E[}Jƙ�,���N��Dw�����ox
7����L�ucX���]rxvg+́�i�e�<��V�'��p�0+��{��1[
#��ު_�ּ;Ⱦs����b�|�y97pO@�{)i��t�K1y�=�U�G+�FzrHpk*�!�#J���_�f�"�$C�s��A	�����'�-S ^|tK=Z��6M`L�&�|��Xln^s�2<x<@!�"��|m�>e�
k*9�Z��T4��m���b�H�p�U)�B鏕7=\Ʀ�2}) ���� ��՚���nG�K�	��^�ܲDPJ�[��W��\�r��w�L�0�Ƥ��u��J�G�/G���\��=��'�ά��RQpnmC�� ���������R'��hIt�ϣ���`q��4�j�W5�UM�n�(�Iһ�(U,��i�,�?L�2g�Z���Gt�
}��z �)�Y�ʿG��ct)���ϔ1�>�e&0�x@�V�#S��PD��b��
�����g�)P5�� �:67����8�F�#Nq���hy��X�w�c�����
d[C�	Ň�d}��;Z�Ea��W�5 ����G:<�e*s�Zv8+��r�pǞid�E��?�v���Ma`4��տ�2ӏxw}���НS�x�N�K������d'l|��T3Ǭ��獖���;h�� ��¨��z�Aix�#����ŀ����;�k�k��ާ[�(qZ1�qK�d��xŗ�Q��vz>��#�oʵ�e����;����?��R��1 xo77�nn4*6,�%�g�&L���ׂ9��� �^Yn}Aj���hDX�/c�y��߲8D�m#F�=hi��0{ ܚ$��3-����d�;	��6��d����=�tfY/7_�mk-
ˤOF}R����f<d�Q��� ���h�s`l�������Zy��3&m馛7���>^��UdwD��9\�
����I8��CU�\�3A���U*�d��@�:��nAt��<�}��$-Ev��u�>a+�k�TZ�!du�e���}�v�DfaR��.�$>3P:��W��Y7ѡ�@T�tQ��κ.�w �
a)��EL�4#�N;����nÚ�df�&J>#*?R�ƢG@�f�D_b�@pv�^�}�U��tQ$�tur��]�5|ʐ�Қ��#G��[]�D8��#?ڶC~�AJ�Fe����o��N{!�0t�5��u"&� HoiæG�P�x��WD�wP������0Ŵ�M���'\��J��:3[��*淒��o%��3g����
��M�}Dh�0-���GŐ�i�ӽ2��y�������Le��9*���5�j��V)e\l@��Q����k��k.kq�ZL~� �ףY��Je�ː�N�k^(�4@F)��SX��G�N��]<ׯ&p��wu�C�?�[_�u�F�c��dg-(ߊ>5����J�%Dpa~�L����7��92���������E�nۤ�Ŷ��98Dɘ�v?�6�J�6��|���
9��wJ�B\e8�s��_tlQ�u4����{6�*品���Ry�~k��Xď��_���0�'sV���=g!����n��[!2���| ��1�GE�6!�;�Y����aK��?�݌}JO'���ѿ��	�l`Qq;�rR�tg��v=(Q��\��#H����C��O��h$�4��dY|�0��c�E�ظA����������f+N�ʮϏ@}�р<�Zʢ��5���x�?�ĉ�E��>A�<s>[��]+W�:�[D(h��'�=�t�N1\N=;�	t��W2lؑ���
cj6��'��DDq�~�g"��N�xJgX 19K��[�����e%"@D����3}dY2���OTc�N��Z���\�t��	k�^(n���_M�R_ �4���������}�yEbN�p2򡒴w���F(��bV�cP��g��-���Z�9�9�F��)����d: �Jm�"0kE!5��Yg�.�U���lVn޼@�+��X�%�1�Wf�ٵC���_90Sͣ�ҡw��;�.�O��֕� �H�wJ��{>�¡z����eTx�1�>8��m�ʊ2@�52r�8��/1w��Z�'�[L����ُc�Ȓ�x[�lv 0��ꑘ��;�4O��"0��Ӭd7��AR�{0��*.y��x�F��߀�Ug�}�<Ms'�T�vW�P|PֺZ���U��
�RR�Z�`�\����F!S�L}�����5<�S�iz|��g=P�@֓��9�8���D�Ԓ�dZ�����=	����j	tC�ǧT�Թ�+��LͲ(_�F
���ɐHE����v��a��B�oy�@T��p�{�������`����y��b����貎r4���c��usM����[7��./ �Ʀ�;g�����0����'�^���]s�&1U<�0C����v;����@&#�Y杅�܇��Tȧ[���s}�vaUS�Έ�s��Q�F�.=g�D�_��r΀�ikvH�>p��˓N�]�Yf������d!����ʶ�=w��<a,|�O�[��zc�[����G��<: �m���B��|�"�_�U&sZ�k�� w��5j�mߗwC����c������!c~�A��|����)ڗ�P�iy�2�ǯ�PjM����Y�l+��O�r:S��"����ח�&�d����������y���d� ����xd��3�R��bx��?x��]�����������8��=�f}���۟KH� ������"[��𺲼Ջ\�Hh�ކUF(��`�B�]�$�Qz�$�0J�֬�%x��C�n$^A��{[���u�����I)X8���O9Z���|�?(�$���+����M09=�������L���:�r���?�$%�ǽ�����r}�@E����n��Z2A�1����ʿ\�5K�{aT�X.��p����;*������Ajq�w�g���ϠYTPV��i/��N���m��Ŗ��� �I��7!,��g6m.·�W�(h��^~|p:�E\�1�w�����&J"D�B�����6�pb��_9�ۦ�$��s(�q�J��Ea��nv�)4	l����I6��jp1�lfE���sv���H��'_�v_��̑f�����g��GM�� )�ݶ��!�E���R1[��(���>4��Ǻ��l?�'���%z�t�%P@�U睙��}��-�,��+%0�[Ow��KXn�'=�>��V��)����豰���$Ϙ0�b�6	�O�JH��)�P�0v՞��Z��>��J2Q���"'����;��EL>���Yv��ͮ���͚���O��� U�ڊspY77���>���|d�h���)I����B �*8�r��~���N%�Pfu���m�/={v�w� vɅ���W�-wTT����R� �R��wi�hv #�!&vߊ_|�$k�/ޗ���$5��5�"��g�t�Z��*r����3�I XJ2� Y�����K��X7N�r=Q�m�lrX�C56���К�~�@�^<������e��d�0��S�}�~�4Q�AW�H�S�"�L���磌���XЃ
������'$��q�M�
k*��`�QB��F��Y/m1�_��E^�n��_��˗��'�϶�����uv� r�&�uν������-s���a����k%���s���x�����aDOL�����H�vxzy�-ЗI�+�JW��ɑ�B{�@�j�k��sЮX�~�+󍿸��H�5��1gZ�b��0+���$���g���c�� !���৴h��Q�5&��M��8�}/濋rmڦM:.|!C���O�-�N�`�9��>@��_���@5�X04�W=���p�'�ٙA2�oFRqs��x�WFĔh���宰�ʀYf�R�_��Rl��t�\Y�3?�g*���~���ܬ�h�z:�㒓3�Z>PE��]S!�7�Ap_D�P��\�n���a?հGD���[�I�}l���fQ%
���:�;DL�}/��ͭ?mm;#��Ѱѭe�a8|\�I�G"�B/��D�+���y���3ҬԙU{��ޖm��z�8zE8��q���@��L6�M�§�G7� �0��ɛ��<�84��C��47\���S�Cs
G&��K?�9f��E�m��7~��	�S�_4���SN�T��M��� �HH�eBe֫o���wj�xi�M�����B/<La=��A2D���ь�%����72��Ď���ڕ�������磥"^�z���O�&,��Z�A�`v���P�G.Kz��=�&>'�a��Jh����H��.-w�L��Ԡ���k�9U���6
�w��vt��B�� �;�4��k�� �n�t$u��rM��c��*j9�l�mQF @�J���z<�>��y��GQH�J��FCf������c#������}x	e��GY���z�'� E$��w8�&9D�<�����K9��U:�;)��g��J�Nؤ..�B�4>�/�wށ�{�|�lp�9��sԨ��D����s[gꟹ��a�$,|,X궶~鱤q������h���2�E�e�\�GE�BfeE��b����A�ۙu�C�
�R�@n��:���l��2�4�5��dמ��E\���н���D���i:�ץ�;���;���T�����?x�U��O�ky�^Hܽ�`&_{TȔ28K�ѽߥG��f��5Z"���v�*��sq�IC����{�I9�V��Ǒ^��m!hD\�QY8����3z�gi��^��$����AK��	6ӳI*��m9U>)HY�q&��x��V��lG��,B|7��W����2	"Z]W�Mr�J("|[�#��V�w~�QU���r!���Ʈ협��% r���_}�h��{�_�?��a� }��0��olƲ���A��U��}m��4�0D��J,��P��T�N��t���
��
x�nJ�W`��e�3CC��[�l�i��=x^0��p��nt˒�:lv���/��g�aP㥵کÜ�8kP�[V~X��;��M�����y2�q���'vx"�vw�����A5��!�nM0L�1�[���@�`S��-Pq���Rx��2���'�q5�!��u:$/ʍ��x����p��۷,�Y���c�]�XW3�q1��>W��C�V��蘾�����1�}�0��-�v���W�wP���A�]PI�X)�uFQ�I��$�EPPCB��;zBa �Q��A��2Y������I7�6Z��mdx�{�VV�P��F�`�4��QQF�_�.[��w��`�e�Ac�߁*Ο���='?����L"ϰ$<7��a���*�R�0�]�ּ��<��/�~�D;A�=�̩�(ռ�[ʪ�Κ#fHt�2��aQ��S���ǳZV�=�O12�^��.MI?i]�^%��{@�ٌ=�f9J�uӧ�e�&)�(�����Kx�&�Rm������m�mm�Bx�3�!rX�&�~�l���_ �>�h��"~�G�a>b�2ay���g��DIddx0�E�m���c�M��&��psT�o��[$�\�S�jÛ�4�[��أM�:ռ֏��Q��?Q"K��LhP3����k�3��5G�Tp�y�g�/��T�jI=��;�r�c��#{�������nM`,�����R9����yu� ��B'�魳���|Ɲ���얿�{x&�(T�:���".G��D��߲�Ĥ3�%P�v<K�gVP4��K���Rף�ԕ)켆�q��1��#2�:���Ѓ���9����G ��,�����&�d�,�`E����ʠ8�l|G���ss�n;3�(�ӻ���癇��tZ�8eX߳8�@��A�>��6f���2y�oVA�2�i(w��4�CI��M��l"�/?�Ȗ�ē��BQ%:'̮dE6o�;1������mRn�":4}�e$����K�X5�I/Z��;�Ie���4�a7Ǿ=���k�o����@�ἱ��Ro��Jks�����9}�%�Q���xGq��CE�0- �OD�Y��	���F��<MוNx%����)�6��<�;w4�S�⿝.W߶�঒s����B��ND�,2� ���l�`��O>ϼ�t�{H�"�}���E�!ma��%�	�����c[-�"DM;C2���î�,���K�FG����H�z�� 0Iƚ���O`��6�G����C�u	WUq���w����>/�Z�cُ�$�m�0��:bʇ�g�X����G�x��iEF��C��'(�g�,Fڦ
}���7���>kH�B�D�:���X_V*akt�P���t=�1ԉC�\ޮ��\�s��k�r�D���ze�����+��U\������z�w��ό�d��C~:�d$����@�e��1�`� ��v��A��-�n"�;�WO��W��9�cФ�R�t{��O�b,n�18�`���R
��,4IB��C��׳+���������&ۓ���P�+^1�-v�i�T�pۂ,Rs�0�RGp��6�U茉���h%����t����}��[���0H�2.��;"A��{#A���F�ܠͿ#'�6�6��~QCso���d�X�N��*����u�/}h��4�-9Pt#@�q��b�'�8q�+g^��m��BXj��r�@D�|��4��4��N��������������ش:B��y�~��c�� ����eo�T�Jx���o�^��h���R��?Z�I�*�toKe���%0+��C��3�������3!�*R�2���	j���d`U��=����u#Ő�ך� �-6J�X�iް�8��=fl��yX:�
��#���/n��B�Չ)����	RZ���ȉX7��{w�����"�[䰠���lI�h�(Z
�K`a3�Ξ�ri�ǣ�VO�Nl�ؾ+ɘb�M�3�EpVS��	{u(_\+���׷�����d�J�s�����/�A��ɲ%aCyD��
M��
��:�=��蹨4�B����ឬ�G�|b}�H��V�z$���i�@��vRL�5N*>�UcM[��R{^��Z�ͨwFA٢���8�W��h�Q%)g�)��ֈWD߹�ǃ��}�8�����uog�X�*ļqF|�*�q�= �g���}K��"�c�Z��9V�?��J�o����� �n1��@nr��)r#~ܬ=���"����v��I�o!�l��,�i�4y�p���U�z����IR3w&o�t�@�6@B;�4��M�mʵ�������(F�=� 󛥯c�¢���ȍ7IW���[i4M�Z_=�tn�X�wl߽���1��ݥ��
e��;\��pve�ݲ�܅!�L��⽾�MmR�q���G@ls��@�B@����K:�J%8�]p�=Zr�ĝ� �~m��d����w&���q�y���$�P�O�c��"뤴���`vOi�G���&�C���hkf����<g?&PkY�����:}�):ջׇ�E?��x*�>	b�[唾ڻlv�ål���g���G8�+ɚn{�2��>±��Ќ��)�v�'�_\H�4��������~���k��yK�IK`�Qg��e�|���$����в������T�Q��ih��=wǾFo$�\�a�9͓�qց�f�Z��v�v&����0n5��Q��<6�j��O	>Z:V�^�q���H�r���L��2�j�. %1L	�$z(�l�g�u��Qx�lT��>��0�L:w�;�Hё�Q_	��Pd���YK&���a��.�q���ꨲƂ�ڬ[��p[VV�m=�{{����(l�S�����6#+n�H4����/��VL+)�2�\��Gk���:��/lW*E��=�_h�L��Fahp�g�˯����%�X�_hh�8u�`>���gI���]M㋫n3o�ro�4瘧`���:4n�����@>��X�-P�V��yh��w�a�Ӧl�^�ފ'ا4/h��h��E�H+�[N�Q�4��C�3�"��/9.� �X���kb��r�2�g���	�G 0�Gz����rP'gT�&�l�B�_��l�<rh�����_\a��V��B�䮨����E Թ�Α?[��-��3)�w�%Ckj�s�;Qa�yz�d��x(��f��=��#�m5��#$~��f���"u����ph�Ω]�	���jDv>�����=��2\~�g�ml`{���&,�Z'����yR"輄|<�>�ô.x�
�K�av�VHŃǭ����u$8v����XNl�d��x�������7xʟ��9��)�� W��/����η��d`�D ��§W��כ4.��b�S&R�T��l�G�R\��W����M��0kF���xa�� D�FG�� ���zRS�!��1˚h��޼��vm#u]��Cٛ����4��M��v0TH��K<Iiq�,�����#N ��Ĭ���D�r5���Lm��E�^J�(�ֆ+%�0e+��Xw��8��@����3O�O\���/�b�D��&+6^~�A�l��h���5j��Dy�R��C���ۑ���a��@�I��{��7�*�;g��/���iti���:V���W3�i6j�_�K��6au#3�4����.��9+D�#��H�����G�GJ�2G�8{u�Cb�s#�ڝK�=���]�6��o�����%$Iz�V,�W&��W�Uԡ����$��'`�
 xE��_2��n�bmR&���S����NX+(#�N�f횎t9R|��C�~" ����'��(�U\�
"��0@j�5���]/&�\�-�vg��3���ל]�.X�������d,G���@n��m�H���Y��#�>T,�����Ʉ��!���A/�ϑ��W�ܟ6��c����1ta�j�e"�bG���?���i�T����8&�����FX�	��B�͒����~�EME��t_�6іsr��B�Mh�����hp�6ŢuU��Ls�D��d.����N�=�iǊ?����|GG�P�+1��Tܧ�\���|g��3�¢�o�ɦ�o ��2�o��G�|(�$���5�n���F5j���"��y�.��YX��7s�ޝ~^���Im�U�rF�H���9��txIWs%*`�\���Mh=���� <�<������e�e��@%�C�J::�\w���`ȋ��>�FQ���e��gYe${/�T��<02��[����n�v-[� ���Aht��6��P�4O�l��P�%�����D��t#��jT^䢅Q��)|I&���3.�{1Z��]X�C:h	"���@M_�evm"f���%"�RОY]O�Kg����2�R��$�~dv3Q�o�"�N�]���L�x��.���:fV�3��FJ�3%�߭5v����L����/�� �P�����w"DI�FԐ~z�Yy�Ȟ��Ek�.�3��;��A4�׾v�0�+#�
D��-�z��u\�s��K��?튏!�ioO�����/>G��aB��b5�";��`Z�5���w(��~|~�1U�~����]_O�5W�Ӵ�������<���:;�m�*�qGk��7��B@
�&�e�y
�?#�4O�z���V�)CϒaB�΁<�����0kq!i�M~�i�R�GH{����!�D���������ӯ2�E��H�;���Fm��$�+x�l�/豗i�m^����(�ど�El��`�䉷����e߂��}�V�o�+f ��%��G:�+W�}�n���"'��m��]'�#��F BҌl|�f��ƥ � 7S�$�P�L��|oX���FYJ������1)9�1s��J�i	^���q�6� �f��C�T[�gf��%�=�a��<u-x'!�v����!��^��Zd��b��":1+Q���j�>���I|���ѭo�X
L:�ݼZ�-���+�������S��"�W7%�IbEY��bR_�rD�7g�i���}b�2
C���f]�%S�/�S5�]@ֳU��w����Np�u�߯P����W��f����b�9��;���d�a�����
�%�	�� ����\<eK��ьi�f�WI|G{W��X�y�/�VzFa��c0�V��GtŲ��6y�,��O��s�7���?eGtw��U�4=/(����`¾����s���]S���2�O�8�������H�9u⛜A0���~Bj��]nda��>wH��\ה�ن�lwI���%Ӓ��Ǩ��b�&FY9�x�_�̢\"��iࣷ�u7���7����u����ӟ��f�_�ekl3'WĐ;3q㒪���"�?���bCr��N�,7��7�E���~��P�~V�DU��s)U�y�V`��s!��#d�.3�4�I�G�??�+�)N?��&x��;����u�d���8��K|��S��y�����d���_ _���i�����:�M���C
d���4��tB�uB/ m?���D�����t@�3��#���yᱺ�M���&
�ш�.5u	���xh���
��Xu�d�iG�uUI��d��Y�Q�'+1_e=��C���w�(�U�<�'~ԘΖ���4uꢟQF��ےr�� ��Z� ��y��v�\�T���0["�������9n�K��S_���S�)�v+<M4}h�Nv�2ٹL��~���m7�"D��ڱ�<���]<Y�EmU��%�	Z�\���uWG�O.|@���j�T4����ᡍ��^�~vպ�}&To��ٛΆ�y�-}�ni�0�U6X�V+�Aa'-�\p(�/�H�w�Ǭ_��%Ql��-՛�Z��q�+���a�l���o"��9U�nf*V�i��+���I�QJ�*(�ҟ*�h�v��Y��YV�Fj7�Q���@Z�SS9b6yE8�0���|Ow�Qρ���ֵ��x�i����˰���}E\�����z�΋]	���7| e}gx���-��������@Pfu���@D��8P3
qtKծ$�������v����V
�D!��ޫ3I���=KP����=��)�� �o���}�����!p�u�E	�����S��ؔ���;rz!F����9Rt��V
# �wp]α7����WT����3�b�M�$'���#1?>����Fe�E��������+O��m�~l�zJ�\���T{�J3gm�&�#]{�	�O`�k�fƄ1��<EhK߮�,Ņv�^o��0����P��Q-����Գ�yǋ�������G��y
G�]�Z�l {�����D�>�S�Í�?�����zUM�	��,(k�ip@FW�1��x:��D�]?��|���\V�$ޠ��uB�OM�h� N���%k���9j���'��\�cЍ^�k�sQ��7���@"23L�a��+��^�
0�@@'��0�'x/;�(_��HHH�Ŷ�0�(�#m��ž���H2�G���n�R��i�(Du�?��a-����0��џ�.�t G��H۪Ց�>�=��6?B%ʸ�zR���U������U�K�x���C}��.Sz�3�&��,������Ƭ�;G'���&w�wz���<�'�15us.8mj&�ì�J�P�T�����M��/v�7a�Vcr�>L�7����b����VD�t]���t.�f�6��yr� ��r��P���Xp가������Y���S~=�s���߃����z(�3Q�X�J�Z8����V�|�����.��*H@I���^|�9�!�C�iԜ�\��/AH����{ᭋ��Zߦbs��".�!����|kǋF�ܠ�\ �>����R��+Vĭz���"�x��ߑ��� Hi���|��vJ���O��V�O��.]�n��܂�	@��Q�g��k�%����(�Ͽ|����̎�;Oޚ�@.�{���v$��b���8���*������G|�(���xm��{ ����|P����/���)+�%���Rz4 ��(�|*�^ԬI%oT��~z=,����{hX�6���x/�8��==�K��Y��]� ���w�#7��$&�[_mŮw��(��K��� ��)�|r��Kd���b�7��+|Z�v�Z'8�XK���ߗ�5iw�:��(
Qƒ��2ְ�
���D04�Ķ̸)�
���_���"s�?�ud<*�K�V0� �-�*H��:q��˅�����db8�����?�A܎�Е��2�����3x/\A�"qiOe�ѻ/a��,��1�E��>�>C:{�K�\����|x(���Ի�M��^$�ڵ3�heD�+Z1�0xvN���Z�ް-�ۑc�r���t�Q6��Dm	i����"���r$0T��<&�q[�H��VM�yj=�Ί1��'����8攌�7��S�p
�jY�?��11v������{�Z�jR%p�
:�[� ����^֚�ʛw�3o�
�ijMx�&�<%�|�F[J݁,�����
�� P`%�2
�wO�8A��%S�1�q�Ed��[0� 0����'#'�1C���x��-������/Ȉ�'��W$�{��(�{1.` |ոD+���D�'^؈k��]��!9˰[T�(U�<_D��|�1G�$<���J ��U�� �+j����H�Ju�$E��_� *Vt,��I�tl(���,��X��HAI���1gG�^9`�������)�*������wN���b0!�+�Ҩt9����$Y���Zo�t����c�XL�S3�g'�o� ;�����(Ȩ���i\��4�'�'�F�}ố��{}'jQۥ�I���j�y�D<����8���O���a(R7PNE�iRP%@��t1�.��ؽ�C�#���q�=�+9�k�o`��k�gi���}aD��<L�A�]�`�G��B��n���҇���ܡ�I+� �cK�cZ-:>�ZJ=14A��;�j68o2��͞��$j4cG'�e��\�C/q��;�0�:hʟ��X7 @�]�>�Jx�M"v��Z3���$gK((����ߩ;��GW���xb��5nũw�hC�C��鴚�h����A_}6�S���&r�ʤd��m J���-�4T����������3�����t�8�s[� �7������'���K{N��'_}C�B�LIS�Ŕ�+�as%o�
h����O
�|��E/ppV����\V2:�U�s�( C.�-`�8���+�jЫ���o֣��M�s�d�a)�F�`��6�K$-|$)p�A�a~��}��_v����a������C���w׳ֶ�$9Ψ�j�~_��2�W+7����|�1+l��<�A�WlY�S����5��[7ך�ԉ�i�N-�ZFh琓\�I���6h���\���#�`�!KQ����B݂P�ǝ4 �xa�wgŤ�-%P0��/>��,t��oq�y�|^�.`�[�r�6�u�X-+�NR���moN%�Q�'q�k���PX�H�1 �@�)����ʂ�a�B���:�5��߾���������(L�aR`�j4}��aOl1��$�mۈ�P_|f2�4h�*c��<��-V߯ �àl|r�m�A��`�#���*�ہ;��H�*�B�?l"Y>o 
����7.]v�n��!��4�s���@D�wA��^r��G�Q%kG�~2>��d�.��z2l� k!Mf#� �S��ٶw@�
��S*��.���7�Ia�T�k�����G`����`��U3r��]�%�U.a�ƨ9�Y!�?�V�'���Q��`K�Sj?�C�G^P7[o#p����k�`��li ֐��!�؏i�2Àm��z����kA�FU�G�ʈ{��FCi�#��܃��m��y;�~6H����{	{���]�o_�	7fֽ%�h�͓nG�@N�����F1�IZ���K�.\�v�ْ�^2s��*n��v\���Ų�6~���ͥ %�#�V�|Î-ɖ_�~��0��;���e)�hC�@:�W�|�� ؆�]���1�䕻�v�ܻ�4ې3*�z�)#�׆��n��2w~�� մ�OfaE�K��%��$��`ߐ
�}-�y�����Vm��ux$C[sº)�{����
 ����a�Ml�C�8E�p�(c�l�A�S�@��_�߷�彊Y�� �l�xZ!m���O����DR"Ә�kG� �'�:f|��0�؀u��|��c��!.�Q�����Ik��q�y��L���so��c���f����Q�4Z�&m�2{�U7u�	����	Q2}o��:{�q�w����ed��Nu��.RBe!?�������@�T�"�KC�R�Ό"����I�*��҈g������`�����JB�yA=z`V�|">P����-�x@�~g?9�)����q<�7i�|�R���a����FP���H�|�3������[c:�0e���|�Gu"P����71��I�Mq!{�D�O�8r!b<(��*�o�k�x�z=�4%�fF�-�Ǐ7��=51�1���Ð��	w�	�O��lM,0�ڐ^��"���6VN����bV� cy��dV�3yM������|��#BT�Eu�.ȕTC�y.�\o�@���o+u瓰&M��W�<`�eq �����]�O$��B�䴭�A}���Y&�ܸ��d!v��Bb�dI�5|^ S�bC�\uB�E��p �s<\)}�a���/�<�t�|���KRD}FH&t7��3B�����`_h�SU�|�o�k��ʖ���'&BN�a��	��y����uB�,�Ɍ&�#��W�i���7�u�Ho����½�zQ��2�2`r^v��˞�A��u̺nV+ �W�	��c ���X�g�#ޛ�|J��e���{d��ߝQ�����6���
'��]VѮ�	큲���2C5�q��k"���/J'ux�����	l�ǲ� K���7��l` 6��~�%*C�ǃI��QrEwU��v���0���;�2���x,l�1�F��Og�w���	�qJ%��If��#0� �4���J����﫯�%y�R��n�%F�+=��O����յoa~�~!
A��K)ص��Q�o��e�*f`w_w��qGy�:pN��P�]�T�˳�'{��X��-,�n�=�U�ب�k�Wt�)e*�A�[�z#�.
�l)-��s1��Y=��c�ڜ�$�5@�ycMp�b��T��o�r$�^v��RS�p��ƌq����ݕ��ĭ�K[}����%�%�'��U�t�S��o��q����-�?X�GN�����}r���ݰ`�Mv4v�K�h������@:~�C��}��[�b�������Eo�F�X�tzMu�����˞9���{^�iH�H��2���P53庢`�]���>���#�������$�t ]�@��ڏ1�Q8��Aw�z��Q��QMB�|\���|p�b�RX����,t���E���b�ߍ�!�ٙ�^U��
S9�yJ���wq9ě�7�Û�E~�oG��:)��R�8I	����_���%�FiOF���P�-���˦<I%���3���5��E���U`������Ri�]�.����G��b�U�(�L������M���ӫ33�3��f[�h�[�^�TP��i~���Պ������?��j�2�3�U}�i��sVj�jJ�,�>4�_���'=�Y�+�D��e����W��Jq�LfQ������kI'Lk� �%��:�`dE^F�8{��E%:&����aE\"��mi�tT.�ܒ�f+���(D�2?Fx>��
�u[l�\J��~g18���)@��:X+H�EM�-T(�v"��^1�v�4lMy��Rݳe���p��z(cES�MHna!�p��*���+5��`���d�z����ɋf�&�P؋)����,S)�罊�"�6Z�B��pq�by���%�MU�N��4�Zjqd�`v+Q%�����t	褦�ދ_�������p�[��U4�����Z�^�@���oo�@#���Kf>(@TE����A��Y�P٪����-�x��x}?�[p�I��s��ya�;�B!*�Ne]�ډ8@Y9ɉ�[gb�Qײ��<�����(�D��Kk��w��v̥9�7G�
Mɫ�I���j۔g@?5��0W���A�P虶��IO��7�r���u҈4_Q;Ӑ��r�d���~�����'\�'e��|�M(r�5x?�W�����^���T[$b�e��D'��I��	�'� s�j��V�sjO\�,���,��"`�3f�����;����4��ӉgQ$Q��\��kҢ�b9��4}�ބ\��
rpc�Q�ŕ�����M�{	
���͆�����:�{k1�޽�{��ݥ�Tq�!/0Bs���;LPS��H�iL�wT���$�_[�.#Xtah�?gq��ۙcpx�u�{��xO�)�ͬ�n鹕󏐟�$���;��+i*w�jG�_��!ٷ��ᘽ=b�ͼ�M��
�~�Lj@YB|Wx�$�!Sv^�^��Sۊ�լZ�U�������2�������Lu���L�SĤNY�Z����ơo)����1N�vm�4��!� ь�޼E�opf ��g�fˣsp�+��UƖ�n:����јY?�L5]���`)�|��U,��w�ɿ�Uzɿ��k- ��M�ou�_�q�6mR6�)�4���M��T1��#�DV*�]584z@Üm痐l�oe���(K��I�r�OL�f�'ک`y�(�#��c�"�V	-�1�w�3�!������S&<�J�1����;j.B�GFo�V!8V�����=2l{�"=ڗ�F.����Z�D����s���{}:^E� �"-���8�CR"lhݛ����rM��0GH�F�|ǭ�#]�+/�/�E�{�0��r�����|�i�����l^�.�2?�K�t�/��(�A������+m=E
Ե��>ƫ�/AQ����� L�~$��]�Y̙GjR��F!S���ܦ�z#B���K�..�ʏ+Q9"4cc�~\U�3/�їj�4��Z-V4^c��/�"k9�i�胜-�l-��*��ade$��A;uT�M(��7�{�q�6Kp|Ci��w�k<�V>���
E�/�/�E�<���s�_��<I$�&Dy��8
��f�M�C^��U���rr[�bk�6�>
�4�~�Zө���c��y�A�!ߜ?���|���*x��A�O����gft�#��`� lH��)���eR@&g��*�,�z��q��Ěa�?�;���υ��>�ߐ8/�Ys3ِ��q�%$c��(L��������*=�0l�B�������hA����4e����������9�9!�������4I+)痑>�_���yƱ�k�+�I��Ľ�kwqp�+R`�ߏ$��a�#��"y���Ci;���*]�N��3�w�����p�PT���ǘjd�8
��~�=�t��Yw�%%�k�tˏa�wW����sㆿ�FV_�C]�&��i}o
 _z��6���R�Ve���lΏ�N?˜�7^?L�$</E�-���`mQ^Py&�X`��p���ߟg�#;X-��^���Ma��9�;x���2�X��?:`Q�N�A����O��X��bǄ�*w�jd��>�R����+>5�Y�����%�7y��fɻ~c��#J�z4���u�TJ$��?����6�3MK�Ps�v��Jˣ:���q H>af <EX�!p�m�����tx�&��T�,1��LrI�-rA���p�D����n�ݒ�5r���r�j����Ѣm������b�~lN�a��]�4<���� ��u�HiX*LH-��7#	&(��%��v����&iX���n8��3�xD$�3�������{1/"_V�������뱼1��ԣ���0~����g�%Q�|q������ Ę�󷤤e���3�����%��V����/�U�W�w8d�FW�d�B�pYV�a�v�eP<��=����ܜ�dg4���D�Z�]�U�#yZ��;!_{�A��'��Qk�ǘ2��*�]��CSCT+����mk�3����a���<�qų����q��$��<ῧ�>���(�ҽec�IRԍ?̣nC	g�-�{;�罷�J�*U����-H��^��E�ؓD.g��+Ej̾]E���'j%�>�Ǣ$��	>�}޲�T]i"�:;���d����=�qG��m�L$��+�t�@�"�3i[M�0+ui.f0K�*���o.��Du	HQp��h@)�*�hK�\q���m��W�A�42��b5e�O���=~��_�ڰYd��17+w���}qaoV%�Sѷ�i�j˱��e�m.z'�!x:��W��u��^�z�1�I\e2�/������y\�>'�D\�㯷#!��S/��e'��o8�*�)`v�; 1�����Q.�/�$>^G֝�Q*��{c5��4LF���,c�s4*�@��
O��O]�nlN��xh��?ʏ��O6u����=�$a�/a��>�F�ɉ�ci#��K�K�h.RR(�'�V��%�V!	�̸���^��Ž�-6�k�Z��(]�������?I����s8d!���q�}��:����k��05)��9i��2��+Q]���V�q���|���_#V]�*㘳ȊJJU�XP�i�α&�FDG�*p�bK���%�t��?��K���T�2++�jCВUEz�K�\�o�e��Udc�����^4����.�v��h��s�K%s"Q��5O~k�7R��:����\��8�0B����m�Fp�3�E�ծ�b'�ى��� θ�1v٫�1�YG9}5A<��#k�v��Tә���p������F����gI�g������~{�!S\b �)Pc��d����V.� �Y�0JI��V�Y۾W�8^Q��t�SZ�+��E/iv�W�U�i<�dp��A{>��C��{GsU�l��|�:�>�����N�|�؀54�Q����W^ȊH��j0s�G���
,�e؁�>��K�y�l�.H���9�r����^�z����a�T�c���S
�FCj�."#s���ډ�Ɍ�����s<�t߻L���a^���#j��[�8���{�{�.��Iw��]�Wk�OI�l�At4���E��ne���+U�+$�	:[�'��>��<{����f��H�P�A��D��#AH�W+P��V���<�Fz�J}·��쀫��yn�Rf��#�e���	P���+�Ҕ���`Ŷ�PXf	�2�F��a/%����GN�p�Ơ��<��?�x�S���	���j~�>O��~#�5,�_;a�����`�.U��%
�b�u����]�/U`f�+І��}'
�d���QT�����F�����_�⳩�R���jq�Ɉ=05��,
��o�vV��m�����l����5<x��!��i�=�t �SI$�M�VOֹ3¿A��}X�G������A��V�=�B�,@��N��X���[?��gmC�KȅŚ�Zx�"`�j�_�#V���h�!H�Q�kǻbp��>�}+i�\#b#�t=��`3����/�4ax��/�fH_
�ڑ9�Dn���J��|��w��d�Y��c@�`��mt]s0d��$�+���i�X�޲�?I����{�5�H��o���)K�@�U$����A&7����� 0�Ȅ63��9�N��5� q���Q���k�vs���W]��ʭ\����1����b%���y怦�
�����
�9_t�8;�+�_�x�K��
N*��������Sر�'ߝ��]�ՎNM�	��a�,�����Ci���9[�Q��0����������fJ�	�}��3֒O��ԟ���[�+?��u���mg�Q��N1?���Zs���{��@�9�ԧ@�M�����ڇ�y�?�VA�P������m�yV�w�� a� �V��f�xЂ�R���O�\��(��(��,��^,�̷��h�[��E�K�_-P�B6��k�,�I�NJ�h.E�fK�\7�O��jO4$hϻ��4��}�AX��0ĵ�NB�7uT�"�����W�Jf��	���v��"����/qF��Ly���P��jGh���R:��Q�m�Y'r�E�S��;+[��y�����Ms�G�`k��d�� �R��o2���XPk�ԋ�fMt̯z��n��t�-��{9^+i�cBiH0,\F��;��Iiz���u�s0�Jm���]��n���� M/�4��P�g�.���QD���8xw��N�\��"���j�-�0ᓂ�����5�̸��5I�${�~�;��N6ƞ�[�D���÷(��T��"�Q�H�����ϼkwگ�/!�ݻ�2ۗjE�LL��Ɲb�:쳛�k�GY��8�X���K�+�:,h���!2��r�)����	���5�H��Ĕ��[g���g���-��f`�*C���{��K������tD󦜛V`ece����EN�J�;ʼ풩�ǈ�>�ޙ��y��2�sҭ��ݢ�v#I�j���ClDYf�l ����v{�|���CI�xg.KP(!�)_��8v�'����DYo��D�@!hg�Kƽ.Ø���d[U[(|&6��4��4އ�)ė�J*�,�&�d1[Jr�{5 u�jhI��l��A�KA��D^}D��S�$��ʎv\S"*Y���z��9��da��eQ�e#����v`�����@=��a�e<��P2��.�����͑�n3`]Kԣ��$K�0|���M��7λT��r4T��9W�yoG��ƞɫ�K�9u�"�������O��[K�٘`}�'��qvn�N���}�L]7��D6��Ul��T[�p�P\�iB�2�$ch�t�����Dg6 ���A_@�"e����R�'l`�w
/up״���~7����A�iB����dk{�� 7�S����T��]lz���x��hG�e1n7A�h/�׃6��q������$s�O@�g�M�pDm�6���*���j�����Y�Z[ţ-�N��}T�P(��P�1����p��
q)���g��;7]��4��/JZ���ϰҪ�3�Pq���P9�%}6���g�*�Ƙ�N�]	r	�O��:2Gdk@elP?�"aH6Ia#*	�$���}d>$m�!�I�s9�2��n��
]J5)N��Q@�&3��h�!�'ơ���Ve^g��<���՚(�W�� (�N?v��=����Ʋ���$�h��\�-���F�}�r�������9�R�T6P�<�5HW��-�0Z�=��`!x*��p�~2Ė%+�Z���O|�>z��э+��ږ�}�D��6o���!d[�kPW\��7F���?��Zo�w�w�`�P��yۭ0/] �N���<.[��cvt$�%W�����C�LĀ8�KUx"댱��!� ֕��oI�����Z8F�me�s@���-��_���SJd��I,�|��� ү1�9rS���A�|�|+8�6!.J��$�e&|����z @(~��-*�a�zR���.�(<���%K�*j'0���v��W��(�IZ�^3~�5����	&�A��lwrN�-Q�������(�.�g�D:�#/z"=7���%��s��A`�������s�wG@��ip/�R�	����2~�ÓO�r�ܕ�g�<�6%�Qj�ݪ�Y�b\Z�*q��'t���s<���ʴ�9�t]�c�]F�OU��:,�k�!*�^>7�R�4�<��zR6�ˏ�A���2^�뜀0HЉ#D��v�q�=h�B&W�	���x��E}F� �gkUL[1�iM�Q�*!�b����b�Վ�<M��%s
)nHa�X�	nq;uٜK �5� ~�,K�HⲐ!��Wk��7��̈́�D��Mn��f;[��v٭+�Euv�>v�a��-ޒ���b�x��+�m[қ�*4�C���X� ����4>��s�#ua�H4{���6%TX�7�����hQΡQ��wu3���Qw����e�V���F�90�a-1�i���R��?�L?~���n�P
��4����b���f$r$���_�n�Ȧ�����GH
��$̙�.s]ժ L�h��IX��`R�.��U���9Z�����Z&����~���,�륊�Q��\�w/xTH�#QYFf��(]�c����a��]��u���s�ն�R����Grh&QhZ�<{��&�3oCM������ݗ��j�Ú?�B`6ghOd����	���m9����6FY���/	�H�!~7+�979��j�o)�����垼4���A���/�����%�?���"�T�t� A�;7����A�/%� +!�A�fi���#�BB�z]N1��H�������IU��M֎�k�x2�]����L5��V1,+�c˥�t\|����_E.�n6�b��Q���e5�����'���ˣ�+>q8g����$V/D9k6khV�ⵋP'�f�C6zc�	?>1s�������7�L�u�	$ �t1�O��Nx�i_�EzI�{����zG�O2 �$�N�D��[ ^le$��d��<T�\���*�����%�މ���`õ��2�{ՇO(�Z.�	����l��E<V3a~8h���K��E����)��aA�1ML��w)��zC�X򗉞+rU*aq��*O�����d0��T��C��r���o�I�"��!�i�s����(H���L5�Qvc+�o�a���b#]�y!�:ߞ㓛۴$�����<�e�������uܙQ�k�U���:ׇƓ�����TX���u� �J�E�8vWX�k��c����l��莣��}�$?�l%�:�&@tT���wA��@̋����ÖVK���%;��0���E]危<t�8Web���		\/��<;Y-���M�����v����~�՜�%�����)�Ak�;�NLo�{i�U���w�"{�1hΘ�)�=�����H����bj���6����F�+Xo%b��C>w��$E��wY�h�T��q��<�9~��z���l�Vf0�V�)v�s�4��$]��+�3�?��`�`�M^�t�C\2�%2Kb��vV�4�*�:)D��7�hk<3�P���.;�*6���P��u�O��*�K��K��厡���r��&gh2�=e����_CW����oؤ�}�䂂���0,�89aiIs��!�&��h�� ��"�5�M��,/��U���T����[�N�Z%{;���˨�__�9G��0��nqe44�H5H�OEfj�Q����A�%��Ŀg���ρ;�O�ũp�E�.��O�s�k�}�	ۡa����2 ���Ř�N���#����C"zuL���~�#����!�|�����0��&] �4N5��v��ɭ�,;�O�l�Dg��{ڦڭ,3d�*4�(��c�ڜUK���}��N6���j'�c�=�ޯ���g,pP=:Jd�@��f���-
|��˦o����g>�` �C�<j`��%bH���3����{�i���8���@4�('���Q˽c�R�4��ρ�_�6Zòw��X�CkX��/��ʘ�لO���Y�����4���%n	oc�iHdV{8YcQ$����M�����6o/�nN<����ʔ�8E?^O��3'��ON���蓬b����;�-�jD+)��j�V��X��%��8�A�5���M������O�?��衺����vAv8��C:V� j�&w�e&_�C��i������ ]���S��
�O��%�e�K��焽�����p5��W���@;�ʈ8�1<�trC�VhGN�W� �����a���y8�Y�6Pv�*uPud�Wp�e�Iʹ�R�]�>�i+��k����ٳ�rף.�-S�B�k
 �l�����TiU�����4�r�.�V+�����C��e(j�q�Ƨ�_�fi�� �sF�B�����-���67��z@���b�gg�!t�"_ӡ`��e�.��>h-����ڊU�����N�7���%,���m��,=!���n*�:��01��ޖVF��̣	=9wU����3���='q�6J�X��H)R]��@A��p��T]��A��2�aZW�ZO��D�;K���_�B�#����Ig�7�w$��:K��؛��m�&61ɼ�X�~`\j�JI�=\�3@�8��>���0�Od֊ۚ��+)9�r�{�?�:����3.4-#�*�j�X�����S,�b���XT<tfTr=af�tN�DE'��tc�l������YN�Ǧ��G_~�]w��!2� ^���h唸x��5�Na��i������������S��3 h��Yr�{�.fd�oV�GD��2��n4��Ʃg9����Y����$�Q�>�m�Ю�DLZ2��Ӥ��ˈ�4PژX�a&2�(�T��7�M���R��5��7�`#�B�a��&�8�P����%x�nM@"DA&	�4�����X�X�`�W���D�VC_�ه�QF8�W�����M�J�'ԡ�����B�5E��g�s�`߅�p����	ƾDAn%܈�e#-Ư�}h��E��[�1�~ߡ��S�26z�-�)d,�: ��b#s�P(LY�jQkc:3�-~����`I��YM蒨�'�qs�8�vv�j���k9�3̾k/�f2��S�!ܶ=�m��f��ɗ/!(�!���hGf�����V��b"�K��<�����߬u���.�N�&��,T�Fo�>�x���������(����,��i��M8�0|[X+}�;"ݚ���o�1��RLm��WS�?C�f�̡3fu�a@�~]43d�!�ɇI���K�A��&h+�¸��+A,��=���Q�P�st��3��e�(|]Ǣ0�dc����l���K����̰���7��"{xv	y�H�R��?u��U�c���h;�u���R!������ ��V����F����fJ�q�o����쫬# �	��vzznT��w��j� �e2��(#Y�gX�����4+V"��	�na�L�lE5��3���g3#q�\��j�W.�\�ђ̱ w�t,Dw�"E�^8���̀�iLD�u����W��B(��i����bl!�uq�R��<�B݀�,�fً�´�V�1�ʱ���ix��-w��bk�{{�t�ª&��������ĮʄƯ	�q��Q�#����X�f��v��X�K̨P��!�6G�#g�8��^�!�9z]���᝽G,�,��\�/�$��oU�w�BO�	֎�+��������Kwͱ�|-U
8��RrsO�=`�y�p]�hIK/on�NI�-��p�������6���=H�	���@�Y�{`�ZΤ	�55(�[�fM�x{�fA"�F_p7�Gi�����Hɺ���Nhp���njF�*��p�i�?���i6��� 3/ ����4K�5��,��Rf���3�#��O6s��W�"{������Q��I�f��Wi��t���w����Z:�z�m��f�/JS��Ec�3C�?�8D����g���!ڛAP�~;Fixa�
���L��qo��܋�.63P��r��)F��8�;0
�㯗��|��V���A�n�Œ��81�➌:*�y�2��J�j����"�x�~�K�K�Ϙ��]��L+��K�
�Ž��$���K��u�ј����A���5�:���p�9�`��!�
S�E�p�Sy�Х�ځ�i���/W���JL��fz��wF��Y]��$@$��@�z0�����{����]���:�P���s	�$}� G�,c|1U��>0�/�@�R6dw���N4��֧	��0h�g��q�#+6n�?I�,}iYx�AA]�9pH���k=	>�+��)����C����u!�:3d���5��6��|�&P"��vs�m�iy��fWKl�)��R�#���K�S�;T4ߌ87u��k�*�4*g�v}�W�̢��[���k(�Y�9�z��Q^S�=�K�k�$��p���/��6V��������^*£~!�AB��a�ZXU�3ͪ�J�\�Aɣ[�;���j�"����C�n�ACh������s�������+@.�8Z��b(�Z���ה��FOY�P:��ʯ)��'���:��M�Q�㷈����2��8�L���UϨY�(W�+8���P؃Ǜ[h}�kɧvG"E8JGvG��?�t���w�Dk�*[��������[�9k� ���>��F�"���	�|�zq�m��B�ڞ9T���J�H-y{��P$�]W;����~��$�m��$�l�p��e"i��3q��j.�����J����G����Q�Eh(`/ا��u6��@���TZqG��`�`��+��nU�J����ǐu��&XkD�#�18�J�M��ʚ�f7"fqפM��j�I��\Y_~m_C$ĉD�����5U�F�m���w�~��/� �m4��\�fd��(��b������.�X���Ft��A�~�#���:i�{�aɞ/-��#��_[�.�kFE�l��NA��!x��B���Y��&�`��;(���,%��tb�fu4t��60�V�K�f�3�>HP~eA�f���/eqW?BF��-�(a�m3�d	�d����}~D�Z�ɺ���g2�+��R�O���A�'�P�R�5}Jf[�Y����E��Ԃ��PM��D�Lk�rDkV!$d��z%��u���T\`��L�$�)�`����t�9��
����Ƚ���7�o_a�q&=�z�QY�l���`�#tê|@Ѝ��a�(6]�Y0b>޴;��/Y�w(	i�a�b'����<��]�-��,_�0�?5��Ĵ�mk�I�>���Y�r������>�*ra�1R��)g��̓�>6�ͲՋ�f����u-6�Ρ��6�����t�Ψx��A���ʁ_hH�d2OS�/�(��pڊ0@�&����\��iMW�N�&+w��!�Q�U '�2dx�ڼ)�*@��p���c�ˑ]t����<`"';�y��rq&9-�v3�<�F�>�t��N�����S���c�˻a��m��V��ʋ�fD��Zr��3T�|��Ў�O�˕M�w��w<plv��$>$�X&�{�2Ϗ���!L��>��́�H�1x��0��B\|��u&Y�b� �etZ����8g�x.�)�,�E��c�9րE������;Q����v�0hA�����3�i1M��ǚQ�i:�ֻ����l�+ �Y�҆|��`9�C�Dq�)(������?@��%��q�_|�����	i��}%g���D��rf~q�T��Gh�6�*�^�lXo��sEP ��q$>a�����H@� �2�QVDO���ن��\�<Y=}�{~K0PA��C�hQz4|���:���>�����m��?!Ӌ2���T,5r�P{p�I?![x�)����X�>���p���p�E�3���߫���KL�1�ͬ�z�D/�1�JQs��]�s�E5�n9�T�|��㿵��2��Z�a�A/�Դ�!��֧*�ʏqF�EP�=���_'\�0�kl}Vo�\�h���3���[���D�v��ۊH~j����
>=��A��n��:4��o ��x��2�IMq�n�Ֆ���.Ȃ%X�����'�k��l��/o�|�8˰d��U�ͭ�GF>�n��X�5�]|	��kԏ�C�%>�w	�|��e*�&uW�.��#�ME���IYT�w�ڷ�JKf*�vM=���W4)z���{�r{��2Wb�
~��9�?
?�0ط�LNG/6��b�!���d!Ι�|�r��m�:>&Z
�h�	$�-.�'j_��j�iby>Q�gA'@ʥLR8j{�A�>.�%c��ܖ�?�S*b����~�Yʦ�G�0�qɒ�8�E�~��&�~�P0��m�`C'�,�cGҐ�Za�/����3h/��^r�R�*k���n|��^��`�q(AՊvQ@D���
�i�6pP�q����U���3��R����Ez!@w7&�Xa��\����YS�#W�1��5i��v�M����j���E���9�F����NVt�~�WO���.�W�����>�>X2�b�_�ͥ;U�fW�D��~�w�e/�а�i͌B{���}�#�h�����I#3�,���U�+}=ݑ��^s芴嶉(�x�h�"+5{y�B� 2�Q�v:��%&�ok��I|��|��u2���/�RP�e�.� �e ���J�W�u���-ӱ�dd��7n}���'aT���J��Pू6�!��	tT�
�4�㘊»9^
M�8��v�����pObpe���yѧ�g���zG�?lh���u�/�X�G�K�1X+h��p�K���:�7k�R��I��'>CT�V)f��$��������Awcm��1X�cS�2�ϺY���R#{�eb�J��y��S�Z��E�i�v`���^�ǭp�^�둡-���n����x�%Ty�:R�$�!���'� U��<dp���-I����'���1��Ծ-�����M����$T��~�o��~��t@4+:��̸оШ=��J�b5a�q�3}��Em-�}��.�h� �7��T�� <�13����o^g�>��zj=]������>��N�Ƚ�c�&Z'�5�]jU�2�nvll���[E�s���B��x��G 2,�J�-��������5����$��V�S �"й�@)�o!���S*t���"p�>D�(��+W��}v��ܞW�N2].b!g<E�jƷ=��Q���F���FLpԳ�-�e(��}���`ꅻ����A�b��~�'�w��1�,�ǈ�A&��g�GBFR�4�K�ӷ�[�t���e��ҕ]�\Z�� ���"�J�R]N`�PG�
����珧Q�L�HbS.WC���Ɔ����;�/�J�ڴ'�=_vFG��Ğr�+�����6�Y�Џ�`�\\׳�M�~��+"�f��Ј�r�]S�`�i�.�8�Cv3M`��G�`���>8d�����L�=�0�7�6= Ү��S`e� �@Z.�T�� bae�o�/n�����)�}���m/�OD&A�B,Ξ���:eK��b�0�8Z�pd��)gѶ���_M@���]�'j!���7~��m�~�.�p��΁��_��}w�Jo�0��)Op���@��r�5|��M��?���vút4�rsƉS�m%�c}H��Thٮ�@*M����������ru�~��hG.x,����L�ܐ������lRz������bź�!��������.X)��,�%�`Ap�⸕F(e���hE1/��|�tx��T����8*�K����~1i\���i�7C�^���bD\*�Uk�S @޽6�G!= ���gN�%(��	 ]b��%�u>�"e��?�I{��Zլ�2�5B%;�a���
�(�;_ ����6�5��6�I�����"��ȉHXA[m=m�n���9�m|�[�؜a7�Ъ|Pr�,��MV ��Y?�\�m/���P����T�'aK���ʳ�=����9�}�_ �|�����$zF�j;��iO��аa�n])�0�c�wF#���(����!����|&�=�<�p�s�]�%I����c�cr���#70M����=wP�q�3c�j�D�W���P�"2�__�,�a2��,d2	!$�_�p���s�+�C�iK��Ő�{+i;4��^(���lJm�~c��P*d\�Ð���ߡ���*N����7�2I�(���5z8(�H/R�'�+A��^��a��b���P/��+-Z'5A�,P���|RJ���}:%���z����$־:�Z�Ȱmj�����P���|��$8)y�;�t#H�#=��PVj|��X��d8�!�ݓ�S/v��
afڑ7N��kΝK���q9]�jZ�V2����Sm���`�=���� I�pě>�����.��f�8�dv���i�Izs�H'QX���Zz���t�!���]ol�ھ�B�3�kcNl����a�s��^���}����NM�IGy��o����L+��/�	]��sn���Y�O�7�WbP���վ�7J�����z�g���/�7�(�u��B#J1>	�J��n�e�A,�FC�嵾e�Gno��4�����D
X�A$(&�x�F�I�n����ѡ�R��a�eǢ}<���;t9���X0���,r��%���^p�xI�J:�l�Z�p8�miuH@��N)�(��� j�y������)���	���΂���d�8�ve\���4�1#����C�r���9,<F�l.I�/ ����,r�n�Ś@8��pL����o���h�}����`�3�;��供��J��+��e_�y޿��t9H��@��L�E�wAE
��C�?�N~��z-~�]�dv���'��༞����2t@��dU)��U�J�K@tP`��LK��?��z���$�D�ƸȀ��9�a{�[�K��4��䝍"�ӏ��po*+���7"28�t�\C�m:Iv�	�7�W×�g{ X�Wގ��mm(=/��0*���7h�v��	vC2�V0��:�Oa�ޱ��	�r|��_���9����Y3@lfJ؍1f+T͟j�g/3����m�F �'yYc��%���6�C���%(��ktE�av��R�R�(k,�_��]�x��?��_<�u��a�;�*/a�<����VA��ԳܓL�&ԭƤe���XFT�Jn�7
�@�'C�*M��q:���~͈��DQ,��h4�Bs�D���\1�b�P<��.�8j��ajb���{gAs��2Bg,{$�Qo�u�(DW���l4��ϗ��.�P�-����#֏������s�,�����VR��j.� ��t�޳@	�Q5�ݻ�G`@)x"���Z⒫��2����< n����Y�����Km�h�.�P�`ܘ��;�?]�f�{�2w��ʮ���ئ蛼��tl�F�|Ɣ��%7��-lA�x�Q�J�'Pa��ۄٰ�|.&.|X�ԞIP(drE]���͔3IYg�E��H5��2�a������f|v��y !���|#
;�h�m
0_y/���	�c�k�u��@��(�j7� ���h�N[D�o�9G;�M`��:�A&쒖'�>'&�^ ���CJ��+lV���L9�u�c�X�(
ui�/KG*G��l�����3��}}�����p�F�Sop�sQ`v���<����4\>�N�vn)P�Ħ5k�jl�Ngߨwy&�n�ȿ��S�Nlr0�d����e�6�����G�E!|,��3�z�`k^Ud_.c��6���M8Yn�@X�� ڂ��p��u���r�C"�>����Y��[=��χ?�7/����rU��j�����O���b�R�K8�4��JFL��M�"���Y3�k�_���+@3����KM�K".��8m
.��Ƭ[Yq�m�+��x9�����ԋ������dF(a�� E�-T�hO	������E��'��
İ�9������}'
�^��+ٯs��s_���3�V���f�����Tpz�������R�eYB�3�wظ'�Ѻ���H��BZK������ h���.��K^��@=�W�v�
l�^��I�\�<�p{���:Ifo�'޿N�SnN����!ej%��Ħ�i�e���*i��̬�����'g�>@U��+.N��l�U3��G��!j3)m{n����Uř�%�9�!�|��	*���E��讦|�M���4�u��!�:9���o��ӭVhG_Rd>ӏ%��{}	`�)-��ϐ<�B�\cq��Et�3���.k���'I��w�V"a�"�MϊE���+1��u��})9S��g6��5FgW:>w�j��
�+���a�bw�I�b�.��LR��W�WC���^ʤb8Y����}J0#�����)�J�Ƙa�������tK��#����F#ڶ�
�&����i>��Ɓ���g����'+���l>��}Z%j��6J8����jar��;�r2�ꟂU�&�qw:�^�-�K�,�:��9fU�|�PI��C[�T|K�uVP�'�����?�f#�*PBg�۔}
(
�����^�v��c�M�fvܥ{��K���������_�C��|�P�ca9؜ε2"tMp� � g0��$_��,D楒D0p|���N $Nb��9�g1�%ē��xb6�u&�cFQf������"o*yXl���k��Կ,�|��ݢ�N���ط0�����H�GXd�,7u2���M;^N���ځ�㥴�����Az�D3]��?5�G����1��W I6�+(�ϣ�2��|@W��x=RM�j3���T8 ���d��f�3u9��A����%=zZ�@ko�4�P�A}uMש��W`�3����/��I�y��@! �I,��9���%3%���>8�)Z­��}�A�1��-��߃<�R�m��~V�n���͌Mi�] d�W��VǤv�zi�g���ʷ�(*j�÷[a�	~�L����+3}���^�ꐡ�Ϧ�4�-�f��+����O������;-���{�X�g\9C��^� r��e�9�b^�T#$ו���U֒�G�WP�V<��T_�Y��}����;��h�$���[ە�<݁�>r�&-���������"K����~�o	���(��M;�)ߠE4?�m�\>A�\v���/��{��l�蔾AެI�z�����B_z&5�����N��r��1h�>%�xϺ�8F�_}^��0�e�����[�K�:�!�}�D=��&y�$����J��)݉�4Cҁ�ר I2���#����/A�&y)�g��=F/w+� ��x�~�� A��4'?l��UG0UX�N�<�"��"\JE_JK�$D'�3��2�E$~9"T�VK�g(�࢓��\ �p�׵�uJ;}>��`�I훙�[_Q�=�α���Z����QY�F�-Ϟ�g&}��tl
��K��*G.l�*��/�E�=x�6���k��g�e+���'�W�y4>��������!���l親^h�Zi�S����N����}�S'2�I���I�"dD�SQ>���'�"ѓ⿄W����l���M�ۆz9F~ub�%�b�����=w��W������Vg1�(����G��X4�Q U͑�х-#���6��\;#�'� ��7�l%H��ߙ�[oJ�}Kc0S:�k�s���+<_ʮ�S�|%g	?��r�畈��x:ĚN�̀-�B�*F�KE�d]��eN���--;�=�d���pJ�_��jܷ���#����V�_o%mc��y�h�����/��!�C`����+�]>m������AO��� wh���]��7�?�9� �N���0��79�Y������mj�R��[3"b�N��"Z�t:�o�0a���.kv��*�_`'�:�}���Ϋ�}�i���ː� �3��˻��?hfx��Wsn�$\�� CA�{:�Z��,����C�t�{?-���/Wz�Ou8
R(�z�],�������ON?�n2O4JzyS�L�ؠ<jm�a��������۔o�����'����:�a/�_q��>3Z5b��J���'�?�Z�����ç���Q���פ��l��a�뷨�|7]�&x.�\�U��Ei�4�t����`o��my�.\�K��g6t��������t�W5%��HPC�YjZ��=s������W�#�S�-0S��w���١�Ls��_�"}��ä��J��.���'�]Xj�Mr��9�V� ��BwOs�D^l0J�,�go�F�5�KG��"�x�]`�(A
��W?�m*�'qf(��l�ut�Q�om��-��8J���s���0[z`_�~s�+���8f�����%I}^&�K��vW����u����=��F��f+�����H�&�(���0����l=�p�C`(����PX�4o3�۝Y�{�c&p���uF ���Cd�R�Z�_e]����L���7kf�����p+���@�Q��Ñ;Tc�c���L�)��_8��N+�w[, s�׀�Wg�[k~t��!�&��x�)�#���	� ��D�I�V(�ҍ�3��U�В�!u�I赳� ��U$�:�&_���t/Vj��uV���,,�Q�����-�����؉�H֕�t��#�$ok-��
�$�Jҕ:���BV9x�.[n(l3߻M�#8�B�ڔ[�v��E	�!% ^{�go��y�/�3|�U?����!J@����5[�|6���
D�8E�������E�Ek+����U{��&ങ�ww^fX5%�<˭G��t���Ê�h+"o�V6�������$V�l���31Q�1�׊,�����:����5g'��yu]���|�{��EފE1�ad�#�2I���`��-|-V�[��r/˰醩��2�z�xu !��L�%���d�sh�$E�P(�	�e���H6ƭC����&c^1��p�Xp'���7��t�Eep�S�|�h���?��i2Å�	XLֺa�����o�xƪ��ݾ�%^(Ӭ���d]0&=�Hv��sêu�������U��0��34�8V0��q�mu�ʧ0]��/��q=1!L�]�X#q�7�M�L��V�����5�-�LBvM 4[�w�<�A��Y�]��K��@��37��	�92`u@��i1S;�J�jI���.��)�z��?,�@�Z.̳��l`7���g���_~��E�� �D`�:d��*f7�"J�fR��H	�i�oT/��;�qeCyFv�@<�=>i����R=��46@�iL��̫��J�'��Ì��|�����Te�����~�!��z�o����L���H�X�/�I�t�͒&/��^ST�S��5!D��LFS/Ql��-��e��pcwN e�i�������z���w�C����Pt�ˬ��^��F�t��İ9��]�����/�f��:w�1Z�W�6*͑0F�:����l�� ��z�*�85�-C���]7⬶?�����ƿ���=%(T��qg(���|57�쵌�2��'�ة4�:��<L��FҩAk�`)m
g�| �D��
��l�ң�0�_���E�%]���`њ,�R������ͪ;�F9FM˝:n��.РzXM:�J��߸Z++S��L�Y��ү�ʆϧ�-HU�1�0V�����56�7�A �xj!q���*=��F�'u2HM5yn���} d��4�ؘ="t`ىP­>�R\���2a�O����,د��z]�}�>wy�/�c�Q��ţ�P�M �/��»lz�``��8�K���=����E�w�W/�=b�}n8�\���(�'^��T@Q���o���dEK�yE{	Y����_�T���O�h)�z�:�,Z�?re����`����&� X���+a襃�d�T�VE�npLlC�?��i��x�ƛ�"�����添��ߎg45��<VR%�R�6��GY6.��`������k��d�	`3%� *d��\+�j_��ݶ�F��Ȓ:hM;�}���?zs����K��7����E���{�Y�q�Ԯ�n-��M�1�˖.y��x6G�?׬������N@���M�On{�e�o9�0d��@.9X��#��9�=r�C���ds����VW��T�dnnG�uX�����4yz����/���mjl� ��-�~��3�s�T�f�9��Э���eETO^sy���su�1f߃t͔��w��.�o�����&t~�x��
?M��Ӧ9G�`�~G��y��J=VwT�����7��E��Yu�9B��$E��'�o��~��F�4'Q{>|3Ҡ�C��M�+��c�eP]Z�E��zEi�ά�T��C�~w[F��.�I�j1��/��O���E�&86�}����ėH��;]=�<͔\�Qv�T�].봜p�u�ΰ�/��mŔm}t�\D��yyѝ�&U�]zQ0�1W�!����rYZ�sí�D�.��-�?�h2��1�䟶ß��õ,���w�.��	���A���~�������-!\��hYP���fk�oʭ�=3g�]~fM3q�5R����an�A�wS�nS�i�OhvT�s�{�=��=��ո�����ā�?����W �ȱ�6�<��[I�ɓw�ivfM�������0�`�"�������Z �˄��
���@h�2#v�/bHo��doP�A�j���;?L.ʑ��eZw�t�*2���k�h���5#bDv[BR����2�v`~=��}�o� o����#�ېABT�ÙG�6Һi7�=�Y�'��Բ�X�?AJ���P�����ߥ/m��b��?Ϯ��8��*����������L]��耸K������C��\�{��<2lY1-Z,���9C��S�۷�2~�n#�Y���ާDr��3�"��
�6��is�E�#�
�g v
�
�t�Y���J��m���t<����=+dZ��K2׃���YN��3�>��X�OB�֢i	mI�!M��c-���9j�2a��I���Dz �g4�5�P�?w�Fj��
�DT.~_<���`�3����ˀ��v�BAl3�����\I���ʖcY�Ðm�u��?���ZhL��]I��~2Hӥ"�T��1�ѣ���Է��ycT��c�Z�K��ͺĺ�4��}R��ζS5�pB�c��G��b�/hNp��P�<��F�8?��V��a`��S�MA�L� �OX��=2| �"�ڹ2$�J���l6�j��%��Q#�%�t"��i��s.A��w�-�,�;��ULܧ��!�
ep���|��t�@�W�-HB+%_;��v�]9I��U�칈��)���w6�dƗF����7�����d'J�G�����npn�\��'t�A���j@t���*K	V ������ :���}���5�d�E�˻�[VP�"?�\؝vb����+��2(��|�{eenO�2���OԺ�Y"������w��X��I�Lwb)':z]r����X���R�l@c)�(���_�|"���Y�|��<�O�b�e�$wK�ѢL���B5�;��a��՘��������Lo�(.���~��nv��P5��:�5\����3ܐ��� 
u}"m�9V��b�2Scv�M��,��,��4��Q�!IS!�'-:(b��g ��^��w��m��ƞ^ ��<1m���Y:з1d��V��亃GI��+q���!��_qP�6k$cl�P�׳�Nyn��V����4�F`n�GqEI��Y??s����9�oy��T�x���-����"ů͏E$O���R�'9�_T�a��@)YWe���	��^N�9����j#�w�v?��q?8Nȯz� _c�cuJ�!fW����|-ɕ��C��Ӏm�� ������IjQt� ������?�Z	�{b*JPyb&�������ϫ{�x�����.5m^�$�J�۞�f05$`�-C9*�1���#�Q/9�l���V���޾!h�Em����q��E�^,8���վ��ǅ�xvx|6�sP���m�G���y)VA�{Ҿ�6����y�
�У�.{��b�ɲ]ZB
�B�숑�܆J�C�3;]j0�]��j��5r!dۭ�����<�S�`���)����R$2��on-�6���j9�⣎\�&=o�v�O+e�Z��D+��R#i�TjPR��X�P'���_��u�<}F�&nNѯ��mH��F+2'��U���!�FrW#CJTc��8�:M�E5��ia�����9)����k:���>q�[AV)����b}LC|6i.g�(W���z��-D���f#m�V=�Q=¬|�0i�;���2��IH��n(���#$�F�cW_�o�GўL�~���[�l��n��"~R�Y&��m��j�p�q]f�g-X�'ôJ�4�27.ƑU\ɮ>�j�/�ܳ��dc��%�2��JZ~�%�>L��0j/R�8�8,�e�� ��( n�aV�E��]�N���l��\W�W����И0�
��6��������oS�"{�4r��B؅�+�%,�IH���~��k�P��Ej��J�s3]�V|��6�m����AM�
}��
a�H��� �6���e>�7A��NI��C\Y����q��~C���_-(ʥ�j�V��Wu��"�H���?-�-=c0^V�q��Ƅf4�b՜	��1 �t����[k�m�v#vw0��Ճ���V棚[�V�bǹqerp�����Q9�7|�[LOؠ!�����b��'��t���O���Q�C�z�k�9 ��kDgi���RF����
�+��u'�����x�8�7i��Yk�WU�mk��gT!�V�<���Ic��۔���GG�t��rL.�v�mI����2c�CQ�d�a�Y$t���;�{�bhw���*��^T�S!ӽ+{l͋�������U(�V��� f�׆����G� k8$�}� aȺd�;p.o���l�R�UXo�fܐ=�"�WMQqtFmKy
<��� ���٠���@���W�\��8����*m�]���ȱ^�R>�9�\�9`�3�Tкpx�g¿���O���L�g����j�?��a��-��t��ri��;�h�#���	t$$���z�\�?%�a]�	P4��w+��Zw��H|-����shL�dpt&!�h--��s���9@nW��Ҧ! 2{���>J��4=c��شSjV�O���,&��H���GY2*�䩏݋A��L3�+�ӱ��ȧPF�q	5
�������<�68��9#�4��8I �d�8���c��Z�f��|�5����K촫\�<�³��c�%m63P�p�
��uX�� �7�uɇ�8�RuX~���g�
c���Bh�K��`�ט�?T�� �މ�|�n�g?�t�W�*���?�.Ԟ��. ^�T������l�4�3c��d��g��-�S�P��_܎�}�)�i��[��k���$w1��m������{���7�V�o�u�I	8.Xy(���6�jE�L8~�,0H��˟Z�hZ�"�n|��P��viHД�FH&�����i�=j�ձ�1����RiHIa7�eÇ�,a{>�Ъ�Q� ���P�R��P��f�S����˹b�����W7�m$�3-P�t��������q@�����6���I!����je'M�dxS����8�T���:�R��ϝ�`�
�O�|���]&x+��������zڰ�HQ�pV@r4�V���r鰖1;��clR	��������
��5��
YK�'��&��/|b�����t�ة��*��,჉A� ��Oy�1��V��2��1�5
�#�0��k��)]�b�~��H�VD,�~�y�K��J�K�\9sF������J,1DKV�P_lȨ�%v[��Kz,J!�	���"��4h ��/D�a�9Ty,F��s��j6��''2
,����
�IU�4�TC�_a��P-�9�x������j
"3@f�M�v�Q�N�D1����!�Ry�JҐ���C�ܑnJ���O�:w"�}�����6[x������@�+�-��W�v���{�@w�y��|�1jdU�{fy�4�۷�*|r����.�qΒ=�����h#��	5�����o�A�]����1�-��Jݘ6'��$n�9�xY�KދW��� �� V�x}�)<(���VР̞��	���� �UW_�w����
0%y>F,c�r�����i�8���f�v{(�,'����c�E�?�b�8AT�m��,c�g6�gdm�K	�tN���h �}H�T������ ���U�/���~�k\J��+KPw�VWOlxo�������H��/^y��v��*���>6�b�[K+�P(���r/����XD>��T�W�@�5��D��%C=����<��8�9�����I�03c���!���3��cq��K�M�n��NؗK�9��J��"��(�����T"ˠ�I��E�'i̝�Gau!@!e6���Zi=ՖΈ��]mjK�+����Wx��k��xuW��D,0U>]#�E��?��0"����S�Z�� �W&�f���9w���N��<ر����	�8��T`���.�6Z�[���mq�dY�Ēe�Bp�)� ��w�@	�F!�!�&t53Ԍ`��V�=�m�Ӝ}O�m���A]s�� ʊI�]cS����	ˮ��gN�_��	쮸�ć�'����m��r2}~V��3�,��Iļ.d߰C�J�C��٧Ը�M��`B�.+���� �M�
T()*OB��z����"����H 4i��`4��58��Ӕ�Q��oOyn �*5ŁL����.��}���߀��v�@9�(���C{�7��P�7�	������Z�c�uM���;b��q���k_;���D�- ;t��{�H橩v-mg��z�y��'.�v��g����Wʨ��a�ٴ�+|W���V�u`�H.Pq��ԔX��8�<ov�l�eV]佥�����9`l�B��!�җ�qܴ�,1Si����%�R���j�؍�4]����X� }/\Ξ~؁�0���6�����4v&_�>����y�� ������T��)��.K3�6��
�/C����7��d.ې7�6^!a��LWp1��� E�"k�8C���1���wM��Q�`(�37V�I6E�͇p��a�Q�k�G|������5軎t0_�5�#��3��!`��ZC��y�KǘڡB'M�̑~V�����O+�3�u�֦�R����q ��c��� ��k�s�ʇ�;2U�ǻ�z�9���%Lj��%0����4cM��R�Dx۾p�9��(�t#
�[�*p�L����n��Iej��Y$�:��Ϋ���U��W��Bk�lKۅ��!�1�2w1G�����)�n��V}���-�0c��v[a�{�=�-��y�f��Y���������Z�j���g`P5\�jW���V^-���{�^�HNY�0�!����}����&8�Eq&@*ye�c�Y~�/��g<T�1zJ��=-�����`ѽ5v��!&�`@Ì���w!ַۡR�A���7���ҹ&�G9]���cy��ͩe~�4�U�D�
��JĨM�]X�s�����L|�/�4֦�v�Ɔ��[� ���x�d�A����w�pcv���-cb#���k��'ŕ1��y9��d�|�o�}l�?����������������P��:�����)he{�B��}TQ���,�%�V�5r"_��=u��(�w9x��2!q3�%guch�7��2��*��#�o�h�;Zr���$?L6 i^#)ޔYKI5w_��ytm�Y0��[n�����W�Si<�������a�\�j����g�Tc倰�d��;��+�[]�Dj�6�	ze>���W��.��1P��&������+���O���'�ۊſ�E}�Z���B��[�;��'#)���Q�A:�~M�A��� �.�~�҈>�����1Z���sq����S'�ˬ��H&'�
����F��'�	��+P u8�qZh麉<��WoF��^��J�����ཙ(���F�o�Fd�ƹA�����g,>�T�g
	�A�.{'�X��2��a�D�*���G�Y�U{��\�v��S_���96�S 5�Jd5fX/���XU�?�r.�����T?���oNin����^#x�7L�v�fs����M���a񨈽^_�֣՟Io7 ��~����ݰ�AH�h�پ��j��e��7�:ifT}dj;-*(��[�+���l�< =zT�3�f���j��?]����o�{c81�*3�&��哓�	�mS��~�{h�������ܨ{_}��h�Z8h�W�-cܼ��-	��#1w����%�����H�eT�s���!ݳ�ې{$��1����&{�.�)�S��yQw�Mzf�A� ��6��B����ޘ��p���?	���+�PA53�.��_f@9	� ��g�$d�X5%�^!�9��p�*��ٴ�w\7�͘����7Wv_�t\��z�l��'@Z�i ��P�T�F��-�j�6R���'�"��}R�$��!�P�P0P.�|�RJ��`8�|��"	�jr �%�a��;[z�<^{�Q>�;�,-�d����w��6,�Q/I��`�x<�JFJ]��Iս�`0m�qE��%!5�jO���>;��G������vE���z���.��qo�>{�z"|��.���|��*:����En�a��N��6z�]��hC�`�Un�/�p����N9c��-h���{u4�j)9�G���A�]�ܧ�>��%�	����/���"�`�ctv����\��
f8�í�,Ksv�қJjY�lgZ���S(�^]�)t\����B���{���Յ�K}�K6:޿~����� 0� X��sġOC����,��}VD�Ϸ��ի�ճ�v'��%�O��W
K5�7A�8x��QX޻$g��V�M�`7��lw8�fQd�V�և�WMlh�ۏ���3�W	�DN��eo������n�LY������ww��bF�=���_�������z�*Ѧ�p`���ꘘ�.ws\;��7�����)��)`t�h�ӆ���Oa|w���j�5uƯ:P��<TQ(����I��L*�{�0ݬn�"t�a�[�Ci�I�>=��%��͙�v5�H�B����E�۬��	�'�ϖ)�^���@�Q^d.�3�f�3���D E�qM���A����LG����������3}���4�&BՕ�<`ٲ�O ���,�Z��G�➇'l�k��������m�Fkæm7^���n��Wi�/�������]tV+�V?@���iXu�9�^�C�NM�5��Jh=���̠i'�(AX�NS����/�>�*�_��O��h@k.��U��3�<Ԍ��E�RG�ΐȏ�&�D�DLRk�8cu�[p३n��\�ݖ�s���m�a� �d\��D�b�Q!���B힗�Ó�t3i���*�\2�����:c��Uۺ�����`��!�To�:7���6JZp�C8LOS b�(czи���(i<=��T�c���Ǡ�}k��S��;�9󇕷w�Ӄ��N�[��E�G7�x��n")a{kq�(�[�c�f14|�k@Y�7����e�up0���^@���P�uY�Q�+�e��)�S����O�3��4s�?����.��h��5�!��浊���\��Z��D�3��	��?✸'�_�$�d�|��]�>S�l��P8��Jp�S�P��Hpho��d��IE�����*�5R�z7��������R��nq�r��V5�NN�2�k��F2�򬲔�鎓�e�nBǇ��?Y����8�nKi8i���ʹ�Z�m!�Ɛ	��5eAkl��`kC���Y$E��/B$+��y����!����?�A�䛦<J�����&��!o[�l@ۘ������d��VM�NѼ9�ě���-<y���|=�ٴ7�0@c�>Q�+��J¾q��t�V��O_Ϯ�ϙUh�{��TR.G�3Q����y�2�'�/���Z:X������j��7���x��Z�qq�"d�q�
�b�n����&�`�&�lj�D>ZPS��yQ3����砆�Iܴ8���3��cWW��yqM�b)��E�;7����~�Ǣ�����ts|i<��ſDt�>�wH�4��,�u�78����z��<8f��<4ܝD>��7\�y��ص�ƞ��߳�l��)�8���·��3G����������yKm���G&����������_{8�������ӥ�P�I/��u�9
�����mB�v�U��mF��ղ���]���{<J8,!�b�w��I�ۘm�qqab����zǙ�`1�nإ�A�K�������	ĸ.V�Z�n��H�s7��f�b�1Q=���+�� \7�Qn�/�C�!���6�6��W  ���ě�m��#=�l�Im'�#G���t��*�,Wf#����O���l��Lֹ]��å����'�wlX2��iZ%��'T3~�|O��]K˄U����>�C�2��x!����99�KQ����6�g�<��,��C �ũ)����l�V�2�o�iOڠEٱ0�28����څ�p]y�ֶ9��y:�X��7l�ـE�������J�w�����W�f:p��p�"�B�gZo�����_a�	:���S����).����S�����}���Bs��z(�©�
+ۈxP�b|t����X	��ɩ�ɉp[n�����p�[�Epk�O�A���s�
v�������Vk��+�C1����� 2^o���� �.���i�C�3w�ϱ��4������ĺI������d�������G��r=�]3e������-Xǃdd\���xf�*�.n#q6���S�㪟b���B�N���?�a�p��F�0-��.L���n_l�qQi�"g����*v�| �����,w������ �ڦ�z����17�"#{�S6��9�.Mf�4y ���ύU`kD�4u��)��f�W��a_���4!�;��TrM�tE/`ї�����<-�}):��
o����dT>�N�'���V�o��9t����J,���Qnb]9�G�{�֠(�L&u�w����k�U �L_u�q��Q	*vPő�)��s0�V�����T�bKN�ϸ�{x1�<ۮ�\��܅���W��
ń�62τO�XM�7�a�(�$&�w<׶,�?��3�m6�H6����_�e�:���gWp�I�/�☽h��H7�[��J��UFKၮݘ��K� ��ZX5H��r�����R��M-r��j8/f�_�UY�+ܣ�qdχ�>���
P��ty�����q�Ա����{�4��*W�uV�G���<�͓�rܙz	KB`e=�5�;�<�+Y7Î�����8��4�w���z�}ݵS	�1���J���xl�N� �r 9.��)�:�]�;��(3cЧ�#�w���i�貕EC/kd&/�c��Q��W�����=;j �g.;����k�.���(�{�DIXE����;��ڞ) 
�T�f��A�{!]�JZd�2F�AF-�>
|�3���e����	��$�����c��^9#�[���
�a����Le�Vc�PR�0�2�Rh�1�DI�UK��'}�x�0����9W��bf\M�)a�,��8�pFk�p	,��6�Yw%7���p�P�]��w���恬Vl��h�gL�Rs�� ���Ł
�L���'�.ס ��W�HO(�H�g�ث1�z��
VeةR��BƉ!�c�e�;��٪��.��HY6"q������@S�C��ii��%��>K�{���ak�w���,�!�M+6�P�E+)����e�˝-���AN��h5�����sz�@�U�u3�����.D��Ն��</&~�6l����Ǵ.a)� �_G��&]Q�xI�-�jg.&����ҧ!j]��O9�­h8[6�}\!��I)Q����z�M��@�z>���F�:��~mh�QJ#1!E�o����w$����o1�~hBp���+��c�-�W��ȃ���S�v\%N����0D�xw�^�K ͦ~��Q����ep�N�מ�	�I��7�[�3�Q�D�R1��g4�p�ª�Y��gԠ�,�04m-�$O\�4zpN��Ic{�~��������G��M����uQ�qg ��oQ��9{�Y�����f�2�FI?g������y�X@�zb&�}S~�j�<*/"��)x�oF��GўS��x]�z����n6ʅ��>ms�k=DA��Z��*ȭ�����f"��UK��eߔ�D��iΆ¢Fs�;s6H{ y��q�~����q��v�ѧ����tP�P;g; N�.�l��	�M<��mPF]ڠ�� ,��9E��D%��ʱ��4 �(��\yo���F E���/rE,o���v�`��梏����P;^����+32<^��]@����m�$ŧ����{2�󱇏\��A�CLDl�k[�kx?����g���!q�{�j+�ߪc�ޯ�7駱�
�ý��^�D�kK��O���@��������!�~�=67��0�{����٪�VY�G��W�(��0�s�#�2��pb�M�x�1P����񶛶p�G&������^���^����1����Lo��w�T3Po��;1��E��ĀWR�R��ԯ��չ�C��#[w����������bm�.LM��Ҕ@��HQ�g�<������
��fz��w�yԸ��D�ן�ԙP�o�#�����6��l�WF������.`ך\?����NLX�6o�c_�(8]�t	i�3��+��D5K�,��	a�9sƎ]�i�->�d��`�By'�EEtkK�{t��K׌�]�Lf:pA�|<��������֎Om2�Br�B] C���b���cO�� SK�C�1��)P�/��Y����Tr�D	*�ZnƉ�s�^��
����L[�C�5J��&eo�U^@͐�_�\qu1S�Co��,*m� �|��ڒ�1-
	U�䂰���j�b�g�~�E@�gr��@�z"�������	=L*�ĩ��ژ�<'`&����E�
�_��7��L^<�o��� �Sה�P �ȷr�|B�%��S_��Ta"B�Qg�F���������pa�e�	6Y���N,���!Ù;���[�=�5q���Jß�
�kB;ex�:�;;G���i[�rv��v�LLa��~��SH�����k�l��i��<�#.�`�,zA W��i�S�p�fN7�V���\>�D�O�I�p���y"@��_�}��؝ϑ*6h�l;�z�p��	�%�P����WkSS�-
�Xڼ�����ʉ�hY��2�����n�P�V,׈�Cg�����΃z�l����[�d��j��oԈ�-|W����#�q"�l��~���C� O��3�38�W����~�Q��.�nҴ�*9�B���q���-)���spv�,�s�Xk��7E�(��:e,�th�DD8�*�k��]�-��y�Q�H����"OH�f7����%����USx����=�TJqd*�O�)�)*Bxw�VB��4aQ��k	 �}���Fڙ���0����:��f)ڂ���}	��|�ڼgH`p}��4�B�8���Bkj�aJ�/�W�2�}���ߵi�AaF�f��Alp�*�r�\["��Ԋ��T�	O��FH /�g^�s'"�����g_ML"�%�����2FK�WOE{Ώ�\��Ȁ�����g�ӱ�2֕�h���m���6ޏ#�^w+m����~����7>E
�	zAS�6"�s_�m�[5S�����t9�x�C��_W����bW>���̺��uuuv�q*��b�t��p$�I����Z`��M®�U�D�;y�Y�j"r�f�!c�!hSa�n pcp�"T�f|W�z=�����%L�@yA,��;�'���Fit�?�HqVڞv���ۨ�����c�Ӆ[Yiq�鎥mw�Y��W��e,�e��,ab�ʆ�������<`j��^��G4h;�z�K0�e_\q������۹���%��j�6n1���M	�P0��4݄���Lcq�ڝ��q�o�}�"���p�p3�QI!�j�2/H�P�t&H\�&��������+6NE��rϢ�ls�����54�Ӓ����@7����z����ņ�v�? �-.����8}��m�L�o�D�d*A�c��E�a�:�b>܏�<�] �����¬Tp�U��#a�v��� =�*�]ߴa'|�3!S�ey6���I?�2�мq�L�e�7b(/�����I��+�$���"�cO���D9�Tt�;R�[jM���¨��|���?��R#��"�0FBZ���u*fx�>�5
!�ྡ�p� �U�S�+��:G�T!k���D�����F�fq����2:�� �,�S�ƟWe�6�Q�l$*fE4����O�7.g�JY�f�2i��W�mپk����T�vҞ[���]��_�V\�[�:Wq�-|����~�>эjE��i�?�PW�$�2�ՙ�V�O"����T(��Ւ6��I���r�kߔ�ô��A�!�n�qU�=�NN�ʮ?;��\��̷%qRc�	؆%m���~��T%'���\�e �(�f}A�B�+���]Ӝ~W2\�����=txL[a8���f���%�?+����ti���1�*�W��*��x~�'��	��zKzB������M��d�6)<�� ���J�k�Ny���`��� ���*�.�liG��(}1
�Y���=m�b-O;p]��2睠����0 �tZM�ߨNp͢���T�L@h���X���T�t�ˮ�T�E��j��\��������5�.��39r����Sۤp�YY�~(
w�H���V���J�ߊ�N��(6\{���^#ϥ�Cn�1O��7Ax������X��%�݌e�X��pZ�y���\d�mC��,�FTA��d/ek�vW��[�U:�!f���Z���>E�_ =o��V�,��V�t�A���3}��d�!t�����)Ꞓ'�Hy�{1Fl���Z� ,�J��k�}}/p�\f^U��$9s��ܔ��|�怐ꖒT9B	�(�uONe�SZ����x���o�vS���z��x�=�3P��i��C��o��1T�����r�:'�b�Vp0Z��!��*YXf��r:-9�x��8~^�҉��6>�-�Ȁ,b7�Ϊ�D�淠9gM%���u��O�$������ �2�`����X���,�q���c1���r����?;v"��������}���;�̊���IY�C����ڢG;]�I�W$�w��1Qo�(K�|������s�+bn8��b�����US�F�*/[�g�Ӹef�U�����4}���m&L�v9l�4�h��wڝ|K����!$_]�W�I�XnA|�W�7�<��濨'(����?�U���t�%m�F������[��u��m\��W�C��pO� irO� O���kXo&���U<�p��Z�,�4��'��	#o�G���)&��t���'�����"�O��Y�^�`2�1��_��/�Zڰ;>?�ft]�E;2�����pr���d_������(���_XԭQ3¦a�r���g��Ss��N��h3���׵ِ}��6��Q�M��������2At~%�>iQ���g��%yK�@R�C�߭�
w�8���S��E;:�vC���������>5�j�Aw��$v������)a������L�#G�lj�c��x�;�Q!�з%������*�h�o+\)OT��<��%�+%���'��&�%B�G�X�L�^�H>�!��q�Kp�̊ǈ\��:W��g+���-� ��F���h��ST|����MÉ~c���}.}f�%J^]���sc�]�g����W?����O���N3c���1M�|�yb�톂)�dH�3b�DQ���ϣSA�X��g5:��������hJ���_V���@^�j�e!I����J���3W�����2�c��*��}!�x�tx.����Q�9x����8P���E����ۃ�C��r{M�%��F�����:b�
�USFVu�u��o�l�.��t�u�;�}4L;*[�%p�K
��\�&���Ձ��-uy܋��I���T�Ƀے��G_�\`��QDl<�=��SZSW3ߛiû z��U��ѳ�#1�����/��8���Iҧb�`�K�u��q?�5@e���"��N��RD,*�V�p�͊�&y�l2@�l�������t��ޮ�M ��:�TVy�X�X�f�l ���O�
�Q/�G�,� ��k'���������(K�I�\�a]�B;��bìI��bq�� ,Z�6p�1't���H��K,��9� ~2[x�����\j�:��V��)�%q[�~4E>:�.�\�>-j:a����E`���9n)�B��I\��J�̈́�'Jh�+�3���z:lֈ�߆��0�����q��f{dJ҈�8�����s�	�0yv8���҅�k28lK%���������B�$�Ӧ�lv���}lNM�Ҙ �T|�k,��,,y��0�"
���#��ƁE�9��LmрoFxG��S��,K��`�zG����Y������>��I�k�uU4$4�:rX��Ł�� �TV(m��tK�v���T��>���̵�Y/d�����8k�E�F��i���;�J�44�6zJ$��� ��T�=�T��w*����VѨ���r+���(��BFYn:RF��B�s��A��V�}U��M���K�خ� ������]���݁�����u�w'ZxD��?����ŉ�7 >.1{�(R��|�/��K0n����d�!K�X�̙>#��$���kƯ)�><�����b�ФT ��M[�,�@�eI���7K�j.�o�q�%C�CL�)47:њ��2��N��E�c*�Iւ��6k�/n����K��KyB:��MA���@��/��\��逾�b9��b���IljP�9�0Sq�$}�gw���CeM#+*�w�-�<�9Ȯ��d�:�^���j�[G�_�3#Ӟ����ݱ��d�A`�H���bu�4�4�8aj�4<�~v����)L slA������u���##�ԡFQ�.$�&�`5�;��CE?�&���~�̨�K3:$*|���pvh/k�V3��g?G���+�;v~�����j#�������2�7��P��E�?�#oy�h�.�sJ�N�)m�z�$5�3�O 4�v�q�y�����#�7��G/C��3����Xʺɠ��ɮ�2��BTW�������7�&�1o������}��`t��O��r� L>N>$r�$Nӧ�����|�͍�UM�v�z|_e��ba����W\3PO.l�5K�����[���>����̃��fz�?j�4�R p�[J1a.Xi�i�]����l�)�H�����`�L�qA�#4��9:�>8r�U���:1��`��a����	M�6��\�u8Yr���|W�	H}RV
'�F���
��4�0���w�-����vf�������i��$������������X&%"��V������I��ۈ�7�+�is��(�$�偂z;8,\�'���I*u5Y"E����(����=4.'�d%���4�v�h�.�@���%�@�zX-�35�Tk��Z�����1�n[{XV����^�?nnMl �R���]<X�s��p��̥�l#	[<t����?&�K��ۘOM.��6��	�/��O�/��e/��6���p���د��1-���S �KS�fi���9��߅z��z�*&�vE|*JT�=��Ᏻ8��P"�훡_����˖�0ؙ������K���2��ת;�Ga:;�-Oγ�.�#��0`�,	Q�|�9��W�L�>����p΀��"����Y�i�ZuV�ɧ�mcXjm�[�i Sj?��8��X/L�������¡n��[���.@|J��}��9BU������Ek��.��C�挛V;�ݮ[�9Gd2�V3�~���e����P}�o�"��2a|_�Z���	HM��
@��V��B�|Sc���1+?><`���N�
*���L.�Ki��"��������(y��J�	�ۃ4�6��N�@�/k����d�)�����.���J��J�qb�a����e]�q�ןb8 ��׈(Pv,/ ��6�������:?��8R�7�eҧx^f�C�\˷�M�`Q<�����~It,+=nN>�s��|�c��2,�xW�����K��i����(������٪7a��nʘ�C��C_t1���` b�i4��� 8T$3��ߺ=i���S
^���"�!B�)�1�s�����S9�aD>;A�F���_�<�=�#2*�g��<��VAW�����p3EN�]w=?�C�&�ܢ��^符�c�WSy���5���0��<��U���?S���K���SB�Ca�R�Y�E����u��~�����wR׭��=I���P`��a��E޷����N+W�=�S�gݣOi�rۯ���d쟮���i�d=?��}q��B)��ﮋ���l�t��0�~�<R�u�lއ�MI��r�@����>�Ѻ�#�E=��K,-�_)ɝ�x����)/%/�d�E�cǅ	���n��[ZQ=I���TqX8c��F1.+f	+��T��S샄��IY r[��e�p�]�9-WT�0y��`��~��s"�7k�f�?:�<���~��Ŧ���q%n�`��10|j$MG��<f��5x6�NsL�/�闰bypdݱ<3O>���yD�'�ɧ^]M��_?�p��2.HR#��|y��r��L�Ｋ����R}c�ʍ�$��[Y�j����~l
���ŷ~��s�&���>�����J##d��m��(Im��->K�J⣨U�}��:Rb�#�j��!mǾ�im��EH��]�� �q�\�h�֒��kغT�C-e4�]=S�X�GjT��{�Q�7z�#�'i�&��ZM�����=|��ڑC�7��s����J�s�����q%�M��&�Wo��� Y�fa�`�,�2���
U�ܜU*�-o1�<֫�q�����T�kC�;�ծ�~;qr�|�	�&3
A��$��uځ����E6,��w=�r������s�J_y]IH@�jC�����|{q*o'g�~ݲLk;d0�]5P[��>5���Ld5���YHL����&����ay"hjN�2�ކy�b�.�� S�����W�j��{��������O����&�e��j���֎�X�61����9V��AI��/Al�'�|D+  ��u(7���=+T�29T5n����,��|-X���m���b49R�<c͕��Ǔ�WW�ӌ�O�i�y�4�|���H��G�o�=�-�N���lb�d#ͤ3��1X[D��/�D�H�Դ�Sv7!��ͯf�b�8� �~4>R���s%I�FCu���q��Sk�ŷ� ��5i��� q!��@�Bc�b���� ������l����ےӘ�mr� ���|	.е1�+���*�mp�q������V]����\Hm%������)z��7�a�n�aOѕ�ڱ�ؠ�eg҄\��z�q��eCU`T�&�Jz ż����k"�j��VIMNa��
��q$wR��&UIO�P���/��:��A���[!'�T�~-z$͂���Q�
�����X��݀��������j��<���CTr:	$��/dN
����t����ܹg祙���oF��ר��N �Kn�.rt��٣?鼵iφ���Hق�D��Og/�]��I[ �V�扸�ѣ
ٟv�Z��(3�����XYI#7'b�$6ư#�^���3p��	O�G�ҋ�1T�&�֏���̨�a��2;�kTް/�%<rМ{t9D�h��`n�JA�F�>yt)5(���b��{B��1��
��j�~��'d7]s��ǖ�:�F����0� �D�?a��8�7R�8kc�(�HtJ����h7k�����*j�w�[�����,=�I�(a�x�.�<4t��>����%ѹR��*e3�((=ȉ��Hl!~�B,�՛0�ǵ�	�޽��l�/�?:��tC`#̋��}x�i�����mv�TRn�{�&$q����ubn��|fL�k�����X�]�d���#��l������u{��Z�MF��$ �t����;��f�i�O7v���i�+�w����8�^��f�~$�J�-��h%f@�ZE� L23`JV&��Pf	ۄ��ǘ�y�Ty��߫;6>�/�'Z�ԫ���@>�m�0���_���څ��Eml���Kև���)D~���7:�]x�oF� d�9A5��i�w`�&�=iX��߾Q��q��KE�80/C�g����;#��I�9�����h�VG�8�ܠ\ ؞�`�@ Gw$�Ҭ���G)T	놈��޽��_�e�t��u����!ԺSgT{40��l��w�mn7������I� ���ev�J�3���![vyc7���E��W���b��3�������݆���j`��H����]��{�ls��~�c�SCZ�]B�ث�:��������j�^²���I�"�[+&
�=V -ʆY�к[�,���t�s�Kg@h܆��9`�ۑ�
���i �rֲ���)�w�`�`��B��۝���0�eHs�3^��\kFg�3ŭ����֊�qk�R~����];����D|�p�G��a��7X!R�!��Qul2���23��#ߦ�[�[*X��:x��Q^�4i�#,׮3���y,@Q�}�p����S��(�yd�{R�c1�G�6��H�GQ��̃����
�Іʱ�G;��X��_�L���I���e�q4:O����f���od?�ƺ�'��T�;�G��I�@��vk�1J:�)?���G�����iTt㘋�8[з�>�E/� �`��9@TX����B`��J:���j����ז,|#�Ò�|~��c]��:�e����'Ĉ߿[��j�\b�T��U����u���uՁ��!�@�R2Hc0�b6��h'ئ��r��'���@B�2�mQ�j���-wu���d���n/lND��WJ2x���p�Vͳ��l;�l��8�rN1x���7�ؘ��Tp<��[���<��;D��j���^ �	�_6)����Y��x"B�汅�}qh\������\�}�podwKu���D�]��W���Jo����Oe�=�о�'�-:Mi�:gS��R�2l�s�Y��/�2�^&)5�&�߄����'�0�q�L�Ϳ3udS �.�*���#��]�����7��/�k���o'��^�.�r��
�獑$9��k�ҞD��*[�>ce/ߜ��B�mD�B�=�ѳg\��2�����HL,7��_��5��<�ZB�v}���0�~u���� .L����oHk��?DpK��������rR�e���	U�qEڬ����@
��q��Z�ZQ�q���[N��Eҋ��^)$��e.U݀\���{�1�s��I>{<hv'��ə�*����N1VE6�w����iҖ-���P�D<��)�:���[wGY��!��K!ݣ��1h������̯zV 6�"
!���l{�\+�u����3��Qͦ�	�UArN>���=�֘�d"�xI�~��+�� �	|@~> B�Kp�A5�k��zf���C����p�$GD����s���X��[����-F^`�s�kHq
$�6hs���8k�ԙ�T= ��������Rم�I���9���B�m�%"z��]q�p�W@1�=s7���/#��7������k8�3�ȫt�]K�
�R����E���d�)no.G�S,�75�!f�&vޥe��=����-�yh��?���֮��	�{n��_(����W�O�{�4ٻ>���Ne��LlD�p�>��K�'����3�/׉��XT9�7���o㩃��5�C	o*�V�j�6�^Z�fF⣫Sv�q!eQ�e��R�{��0V1���5%�x7�X��Y��� ���Ö⍥���!��(�e���pӶg�6(J�[�8(�ޖ�=�3��nO���L퀖wo��IB@��o{�%�_'P�:�*q<�M���\�WŴ]1�j�|
��Ry�2@��Fӯ�\Lb��n�z��;���<�UFׅ��1c�2z���e�v{�O$�2B�E�lN��ߎU�U7�$�R"�����ȷ��H���?O@�N��l�n���VAg,�'I��!�W�:���nڠc{8v�F/���)ЈR��Tђ��yS�IȢ�$P�t�LY)L���)=�.�O�>���=��K ���}sˉŷ�t8<�� lA�]�$�,�.�T�i���n�5�!����������Ğ���kq�7����$�<���^� ���b��ܥ�������-ܦ�<�.�͛�k�z� �f��(����h��$�ݷ��� /L��4�����4�)��"߹�7�&^$�e�E�9�F@D�L��A&b�! ��ҋ�g��e��*9B��v;Ύ�XD;�PH��|�צ��5F�@��g�0�I��~����g�B�>ho���
����N�z98��������#��3VL�bS��!*u��=#G[ȏ����AJ؊�+�����!xs�G�]��oO	$j4���F��&!0M�����c�~�=7�\���VƉ0���Nb�\ty�h�=	O�ꍎ����(��������@��MT#��U���Q�5���:s�;�
+��6Ĝ�|
��"�ԁ�+Ƀh�Q�t��d�gI�Yɟ�&kL%5�`�r�e�l�Eu�A���Ǹ
\U��,b�;�w`�m�X4%���k����3�u��[�s�������v���?
�)Fq�y4���h߿���w�P�^��\3���%�SM9���Z�d�L�]�4v�z��,�3���q��)��ˑ�/3'�'!4����L��j ��N����'\��.�Lf�����e�N�b��'�p�L ǈ��m�Zx�� ����J������|G|m�?xc{��/P�]L��LL���WL��<�Ĳ�?��n��}Ȗ	6}�L��bO�%zB����k�X��Kr���F������ͬ4Bu	~�aH,y��&�K�k�c��f�9%�^Ws�	P\U0('z�����?�6���y���U�}ݏ�t�e�B��L�n�"�=!�q��}Cl΋�������ky̷��H!�쁎֎�b�������Ѣ���$ݺZ��#��+*CX�0p�f��������E�/�Eì�j6�q��G�|S���Dk�P�o�\ �c���9˅޺�s��{Ы����`r;�e�"�h�F���j����н��Y�������"5�9���
�*ӀW�=��cK��UKA���z��G�ϵ��Ǫ�H�^�CJ�ޙ��:L���eQ�>�&�~s��$W��r˥�H�2�m����n�0pn�"�}3�ó�07�8�T�/[�du)"�{0:i;;�5<c�h������ a�!�Z��#4�� ���H�̖�Sr9@�Iz��Ё��*?C/~��w ��i�Y���:��=Ĉ�P��vޠ%~=��TcSqZK���E;?N�x'h��T~wA�M~苅j���Gl���ĉ�5<k\��[��a��Ƒ�V���?8"r֝k����9�VE]�Z���\�	�܀���gL/?�0�ݝ�]V>�7��~{q��6��-zU"�e�$ѓ?��v\�^���L����Yf��y�l���ŢM����rq�Dg�+���m��_�XI�*��:M��<TtH��}����H@�7EmM5��']����T9�a��Vk"����U{��p6���� ��x����BZ���
+����J���~-���0��2�kPi1�}���Ѝ-Q�w����_��D��9w]E�?9��y��L�V;��E*ǁi�� 醗}��/*׺ʗ��n��'��U�����C����A+?4���+��<-�b��	���S�[Y��򝭈�%��1a�~?�R'2H]�%��E��f����Gu;��3 asG8�m6�@����ßk�`PMn �8��8E#h�i�ͻ��:|����Z9+C�/�-0*L��R�Be����H͒���v#��"��`C�==s^�]ߕ���?'�l.�1�&�\ўp^�-��GN�t����=�Sb/����S�ܮ�[a���&�,���,� ���VE��c����
����ąN�.o8�3<����#��NE�Ѱ�?�jB�ngXa�9h�R�����:���BgI��q�g�?gN���!��Sz~�r�<얇ǣ��7��8����9���}�:=Y�Ur���}g:S���D���vd�3:=|�E3zb�+Ҩ֥�.��Q���@$��:�;Wo�����͏L�����:+5e�n�O�~
�����&���|�
����gl[M+����s���߁s�ހ��7]��X�&��~9Ѫ\����,��X'!�}�f~1m����;P��ޮ�+�;n���N�n���_�����4,:��|JY����ӡ&b}~��*6�8�s��Ȼ���v̻n�>����(n�a<୚��N�0~�L+�{�F��μį���%7Ţ_���Zc߁,�f�%�)�c��o�����'Դ�@���ЂI|�M1���ꡑ�߫�����Ic�B��8��'��D����A�,XTb3C�-30�2���e��t�rr�1��l*�D�27�s<15c��2F�x4wqb�b#,���[a����}A��ٲa��%��:3`��$�RK- ���)�.�_���r�a7v�x8����_�eӐQEޒLPfK��W+�ڏzz���ņ�͋�k�OX��VĜM���8eF�7֧����ހSp�Kݱ�Y�0:���FJ<�U1ny
�Lw��>��Vꈏ�ܨ	�ťj��ba���(U۸��Xz�(]��ܧ^�Hʜ����N����	?dzt������2�t��x!�~�����OWy�E�D�����00*�l��߯���?zzZ��	�Jh/�#�:P�7��b���qmMf�М�Z�a���f���s$LtuS�)꣰�\�{N�q�.d�2G��wy�8�+8�곪[+����&#��+�V-kR
��ȾT����I%E�PsG�Mc+�u�fp,Xmy��e�,E��d)D=t���V<��G,O�Wm{W�(���	�T��y���s+�\�)^]��,v�N��=	�zY��ٮ�e��	�o-��+FR���b�^��k�Sg�%Y�n�>;�lӎ�w�bHs�΃�{��	y'Q(�X�M�����.Ф�i��ɧu�8��ͥء�*��DԅZ�'8=r��*�:�b��&pI/��W��Lo�D����M_�+p� F���|�����U�r� ���Q�£u�&����#p�E�p�y bL-�vgB�彰o+Tn���	�\A��(S�n��7���A��+[�V�콱}g���U�`�络K���-�Ff�lvΣe�p^������ej"SK�Q�B�d���.�Z���Ik��	~U��r�C�8�娝�ֽm,��+��$g��02�Z� ]��,�=�7��H��յ�N=Ơn0�]�DwH`�E/3n�}pU Z�b1S�������y+�Y,�H�)��L�n��zJ��;�.*�4�����Y-�P.�8t��u�=mk���ق_�Ƣ�^��.l����wh/{�˱A�����XE/^+y�46us�Z�I�R��9�]`��i�x��\��v�Mh-���#D��zîշj&N_���H��8iK���Ɲ��A������;#>�,�z�#��[z��{\UM��I���#�z�GD�j�5+z�?IiH& ����Ty0���\���~?����ZU�'i�	C\��.�J!έl�0ŝ���WQ�I &J����ڪSy���Ȕe%_t�+a�I3'�`�X�����*4�u'�A���~ZnsʍJ� h.��;3���\G�o��_��]@O*;���ͥ��m� ?�����l�^0�ȝ��f=XD&���g�v�DaAv]�_�g]���؁+��Ľ3��|AT�)�(���5���?�w0��/�YYӠ�C�����.��U�Fh~��#�^���v/N4��4����y��M��?E�avn�,�.��f#b&Q���pF�k<-�Գ����%*񿹬莊QԉL6ˣ��Pl����I_�q�B�o�>���ͭk,�ry6��9���f"��n�Ӣ_c��4$�>��,����a��\oA)��������eK�n�Lv�_����f���ꏸ�#����	�8��W伞8&�
�%�=�V�����8�����C��o�x�Ĳ�>�⿄�Gw��xs���;2����=�gX��4U��x@Q����u+|c���(�N���bLx�ص�֜����t�J��]jSL����j#���)!X�;��'���E,�.d���X�j�w��qM-�=|��*-� �@�|��<�aJо��>����m�+��<:
�{�6�ᖢ ���4R(��x߃������ԕᮭ.��#�gL�<